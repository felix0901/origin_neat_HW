`timescale 1ns/1ns

module gate(
    input a,
    input b,
    output c
);

assign c = a & b;

endmodule


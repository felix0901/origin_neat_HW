
module circ_q_WORD_SZ64_1_DW01_inc_0 ( A, SUM );
  input [63:0] A;
  output [63:0] SUM;

  wire   [63:2] carry;

  HA_X1 U1_1_62 ( .A(A[62]), .B(carry[62]), .CO(carry[63]), .S(SUM[62]) );
  HA_X1 U1_1_61 ( .A(A[61]), .B(carry[61]), .CO(carry[62]), .S(SUM[61]) );
  HA_X1 U1_1_60 ( .A(A[60]), .B(carry[60]), .CO(carry[61]), .S(SUM[60]) );
  HA_X1 U1_1_59 ( .A(A[59]), .B(carry[59]), .CO(carry[60]), .S(SUM[59]) );
  HA_X1 U1_1_58 ( .A(A[58]), .B(carry[58]), .CO(carry[59]), .S(SUM[58]) );
  HA_X1 U1_1_57 ( .A(A[57]), .B(carry[57]), .CO(carry[58]), .S(SUM[57]) );
  HA_X1 U1_1_56 ( .A(A[56]), .B(carry[56]), .CO(carry[57]), .S(SUM[56]) );
  HA_X1 U1_1_55 ( .A(A[55]), .B(carry[55]), .CO(carry[56]), .S(SUM[55]) );
  HA_X1 U1_1_54 ( .A(A[54]), .B(carry[54]), .CO(carry[55]), .S(SUM[54]) );
  HA_X1 U1_1_53 ( .A(A[53]), .B(carry[53]), .CO(carry[54]), .S(SUM[53]) );
  HA_X1 U1_1_52 ( .A(A[52]), .B(carry[52]), .CO(carry[53]), .S(SUM[52]) );
  HA_X1 U1_1_51 ( .A(A[51]), .B(carry[51]), .CO(carry[52]), .S(SUM[51]) );
  HA_X1 U1_1_50 ( .A(A[50]), .B(carry[50]), .CO(carry[51]), .S(SUM[50]) );
  HA_X1 U1_1_49 ( .A(A[49]), .B(carry[49]), .CO(carry[50]), .S(SUM[49]) );
  HA_X1 U1_1_48 ( .A(A[48]), .B(carry[48]), .CO(carry[49]), .S(SUM[48]) );
  HA_X1 U1_1_47 ( .A(A[47]), .B(carry[47]), .CO(carry[48]), .S(SUM[47]) );
  HA_X1 U1_1_46 ( .A(A[46]), .B(carry[46]), .CO(carry[47]), .S(SUM[46]) );
  HA_X1 U1_1_45 ( .A(A[45]), .B(carry[45]), .CO(carry[46]), .S(SUM[45]) );
  HA_X1 U1_1_44 ( .A(A[44]), .B(carry[44]), .CO(carry[45]), .S(SUM[44]) );
  HA_X1 U1_1_43 ( .A(A[43]), .B(carry[43]), .CO(carry[44]), .S(SUM[43]) );
  HA_X1 U1_1_42 ( .A(A[42]), .B(carry[42]), .CO(carry[43]), .S(SUM[42]) );
  HA_X1 U1_1_41 ( .A(A[41]), .B(carry[41]), .CO(carry[42]), .S(SUM[41]) );
  HA_X1 U1_1_40 ( .A(A[40]), .B(carry[40]), .CO(carry[41]), .S(SUM[40]) );
  HA_X1 U1_1_39 ( .A(A[39]), .B(carry[39]), .CO(carry[40]), .S(SUM[39]) );
  HA_X1 U1_1_38 ( .A(A[38]), .B(carry[38]), .CO(carry[39]), .S(SUM[38]) );
  HA_X1 U1_1_37 ( .A(A[37]), .B(carry[37]), .CO(carry[38]), .S(SUM[37]) );
  HA_X1 U1_1_36 ( .A(A[36]), .B(carry[36]), .CO(carry[37]), .S(SUM[36]) );
  HA_X1 U1_1_35 ( .A(A[35]), .B(carry[35]), .CO(carry[36]), .S(SUM[35]) );
  HA_X1 U1_1_34 ( .A(A[34]), .B(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  HA_X1 U1_1_33 ( .A(A[33]), .B(carry[33]), .CO(carry[34]), .S(SUM[33]) );
  HA_X1 U1_1_32 ( .A(A[32]), .B(carry[32]), .CO(carry[33]), .S(SUM[32]) );
  HA_X1 U1_1_31 ( .A(A[31]), .B(carry[31]), .CO(carry[32]), .S(SUM[31]) );
  HA_X1 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A1(carry[63]), .A2(A[63]), .Z(SUM[63]) );
endmodule


module circ_q_WORD_SZ64_1_DW01_inc_1 ( A, SUM );
  input [63:0] A;
  output [63:0] SUM;

  wire   [63:2] carry;

  HA_X1 U1_1_62 ( .A(A[62]), .B(carry[62]), .CO(carry[63]), .S(SUM[62]) );
  HA_X1 U1_1_61 ( .A(A[61]), .B(carry[61]), .CO(carry[62]), .S(SUM[61]) );
  HA_X1 U1_1_60 ( .A(A[60]), .B(carry[60]), .CO(carry[61]), .S(SUM[60]) );
  HA_X1 U1_1_59 ( .A(A[59]), .B(carry[59]), .CO(carry[60]), .S(SUM[59]) );
  HA_X1 U1_1_58 ( .A(A[58]), .B(carry[58]), .CO(carry[59]), .S(SUM[58]) );
  HA_X1 U1_1_57 ( .A(A[57]), .B(carry[57]), .CO(carry[58]), .S(SUM[57]) );
  HA_X1 U1_1_56 ( .A(A[56]), .B(carry[56]), .CO(carry[57]), .S(SUM[56]) );
  HA_X1 U1_1_55 ( .A(A[55]), .B(carry[55]), .CO(carry[56]), .S(SUM[55]) );
  HA_X1 U1_1_54 ( .A(A[54]), .B(carry[54]), .CO(carry[55]), .S(SUM[54]) );
  HA_X1 U1_1_53 ( .A(A[53]), .B(carry[53]), .CO(carry[54]), .S(SUM[53]) );
  HA_X1 U1_1_52 ( .A(A[52]), .B(carry[52]), .CO(carry[53]), .S(SUM[52]) );
  HA_X1 U1_1_51 ( .A(A[51]), .B(carry[51]), .CO(carry[52]), .S(SUM[51]) );
  HA_X1 U1_1_50 ( .A(A[50]), .B(carry[50]), .CO(carry[51]), .S(SUM[50]) );
  HA_X1 U1_1_49 ( .A(A[49]), .B(carry[49]), .CO(carry[50]), .S(SUM[49]) );
  HA_X1 U1_1_48 ( .A(A[48]), .B(carry[48]), .CO(carry[49]), .S(SUM[48]) );
  HA_X1 U1_1_47 ( .A(A[47]), .B(carry[47]), .CO(carry[48]), .S(SUM[47]) );
  HA_X1 U1_1_46 ( .A(A[46]), .B(carry[46]), .CO(carry[47]), .S(SUM[46]) );
  HA_X1 U1_1_45 ( .A(A[45]), .B(carry[45]), .CO(carry[46]), .S(SUM[45]) );
  HA_X1 U1_1_44 ( .A(A[44]), .B(carry[44]), .CO(carry[45]), .S(SUM[44]) );
  HA_X1 U1_1_43 ( .A(A[43]), .B(carry[43]), .CO(carry[44]), .S(SUM[43]) );
  HA_X1 U1_1_42 ( .A(A[42]), .B(carry[42]), .CO(carry[43]), .S(SUM[42]) );
  HA_X1 U1_1_41 ( .A(A[41]), .B(carry[41]), .CO(carry[42]), .S(SUM[41]) );
  HA_X1 U1_1_40 ( .A(A[40]), .B(carry[40]), .CO(carry[41]), .S(SUM[40]) );
  HA_X1 U1_1_39 ( .A(A[39]), .B(carry[39]), .CO(carry[40]), .S(SUM[39]) );
  HA_X1 U1_1_38 ( .A(A[38]), .B(carry[38]), .CO(carry[39]), .S(SUM[38]) );
  HA_X1 U1_1_37 ( .A(A[37]), .B(carry[37]), .CO(carry[38]), .S(SUM[37]) );
  HA_X1 U1_1_36 ( .A(A[36]), .B(carry[36]), .CO(carry[37]), .S(SUM[36]) );
  HA_X1 U1_1_35 ( .A(A[35]), .B(carry[35]), .CO(carry[36]), .S(SUM[35]) );
  HA_X1 U1_1_34 ( .A(A[34]), .B(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  HA_X1 U1_1_33 ( .A(A[33]), .B(carry[33]), .CO(carry[34]), .S(SUM[33]) );
  HA_X1 U1_1_32 ( .A(A[32]), .B(carry[32]), .CO(carry[33]), .S(SUM[32]) );
  HA_X1 U1_1_31 ( .A(A[31]), .B(carry[31]), .CO(carry[32]), .S(SUM[31]) );
  HA_X1 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A1(carry[63]), .A2(A[63]), .Z(SUM[63]) );
endmodule


module circ_q_WORD_SZ64_1 ( clk, rst, rd, wr, full, empty, data_in, data_out
 );
  input [63:0] data_in;
  output [63:0] data_out;
  input clk, rst, rd, wr;
  output full, empty;
  wire   N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192,
         N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280,
         N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291,
         N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302,
         N303, N304, N305, N306, N307, N308, N309, N532, N533, N534, N535,
         N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546,
         N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557,
         N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568,
         N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579,
         N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590,
         N591, N592, N593, N594, N595, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n1336, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736;
  wire   [63:0] nxt_wr_ptr;
  wire   [63:0] nxt_rd_ptr;
  wire   [63:0] rd_ptr;
  wire   [63:0] wr_ptr;
  wire   [127:0] queue;

  DFFSNQ_X1 nxt_wr_ptr_reg_0_ ( .D(n1610), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[0]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_63_ ( .D(n580), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[63]) );
  DFFSNQ_X1 empty_reg ( .D(n1609), .CLK(clk), .SN(1'b1), .Q(empty) );
  DFFSNQ_X1 nxt_rd_ptr_reg_0_ ( .D(n1607), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[0]) );
  DFFSNQ_X1 rd_ptr_reg_0_ ( .D(n1544), .CLK(clk), .SN(1'b1), .Q(rd_ptr[0]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_63_ ( .D(n1608), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[63]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_1_ ( .D(n1606), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[1]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_2_ ( .D(n1605), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[2]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_3_ ( .D(n1604), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[3]) );
  DFFSNQ_X1 rd_ptr_reg_3_ ( .D(n1543), .CLK(clk), .SN(1'b1), .Q(rd_ptr[3]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_4_ ( .D(n1603), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[4]) );
  DFFSNQ_X1 rd_ptr_reg_4_ ( .D(n1542), .CLK(clk), .SN(1'b1), .Q(rd_ptr[4]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_5_ ( .D(n1602), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[5]) );
  DFFSNQ_X1 rd_ptr_reg_5_ ( .D(n1541), .CLK(clk), .SN(1'b1), .Q(rd_ptr[5]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_6_ ( .D(n1601), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[6]) );
  DFFSNQ_X1 rd_ptr_reg_6_ ( .D(n1540), .CLK(clk), .SN(1'b1), .Q(rd_ptr[6]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_7_ ( .D(n1600), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[7]) );
  DFFSNQ_X1 rd_ptr_reg_7_ ( .D(n1539), .CLK(clk), .SN(1'b1), .Q(rd_ptr[7]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_8_ ( .D(n1599), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[8]) );
  DFFSNQ_X1 rd_ptr_reg_8_ ( .D(n1538), .CLK(clk), .SN(1'b1), .Q(rd_ptr[8]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_9_ ( .D(n1598), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[9]) );
  DFFSNQ_X1 rd_ptr_reg_9_ ( .D(n1537), .CLK(clk), .SN(1'b1), .Q(rd_ptr[9]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_10_ ( .D(n1597), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[10]) );
  DFFSNQ_X1 rd_ptr_reg_10_ ( .D(n1536), .CLK(clk), .SN(1'b1), .Q(rd_ptr[10])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_11_ ( .D(n1596), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[11]) );
  DFFSNQ_X1 rd_ptr_reg_11_ ( .D(n1535), .CLK(clk), .SN(1'b1), .Q(rd_ptr[11])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_12_ ( .D(n1595), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[12]) );
  DFFSNQ_X1 rd_ptr_reg_12_ ( .D(n1534), .CLK(clk), .SN(1'b1), .Q(rd_ptr[12])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_13_ ( .D(n1594), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[13]) );
  DFFSNQ_X1 rd_ptr_reg_13_ ( .D(n1533), .CLK(clk), .SN(1'b1), .Q(rd_ptr[13])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_14_ ( .D(n1593), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[14]) );
  DFFSNQ_X1 rd_ptr_reg_14_ ( .D(n1532), .CLK(clk), .SN(1'b1), .Q(rd_ptr[14])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_15_ ( .D(n1592), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[15]) );
  DFFSNQ_X1 rd_ptr_reg_15_ ( .D(n1531), .CLK(clk), .SN(1'b1), .Q(rd_ptr[15])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_16_ ( .D(n1591), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[16]) );
  DFFSNQ_X1 rd_ptr_reg_16_ ( .D(n1530), .CLK(clk), .SN(1'b1), .Q(rd_ptr[16])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_17_ ( .D(n1590), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[17]) );
  DFFSNQ_X1 rd_ptr_reg_17_ ( .D(n1529), .CLK(clk), .SN(1'b1), .Q(rd_ptr[17])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_18_ ( .D(n1589), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[18]) );
  DFFSNQ_X1 rd_ptr_reg_18_ ( .D(n1528), .CLK(clk), .SN(1'b1), .Q(rd_ptr[18])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_19_ ( .D(n1588), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[19]) );
  DFFSNQ_X1 rd_ptr_reg_19_ ( .D(n1527), .CLK(clk), .SN(1'b1), .Q(rd_ptr[19])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_20_ ( .D(n1587), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[20]) );
  DFFSNQ_X1 rd_ptr_reg_20_ ( .D(n1526), .CLK(clk), .SN(1'b1), .Q(rd_ptr[20])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_21_ ( .D(n1586), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[21]) );
  DFFSNQ_X1 rd_ptr_reg_21_ ( .D(n1525), .CLK(clk), .SN(1'b1), .Q(rd_ptr[21])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_22_ ( .D(n1585), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[22]) );
  DFFSNQ_X1 rd_ptr_reg_22_ ( .D(n1524), .CLK(clk), .SN(1'b1), .Q(rd_ptr[22])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_23_ ( .D(n1584), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[23]) );
  DFFSNQ_X1 rd_ptr_reg_23_ ( .D(n1523), .CLK(clk), .SN(1'b1), .Q(rd_ptr[23])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_24_ ( .D(n1583), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[24]) );
  DFFSNQ_X1 rd_ptr_reg_24_ ( .D(n1522), .CLK(clk), .SN(1'b1), .Q(rd_ptr[24])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_25_ ( .D(n1582), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[25]) );
  DFFSNQ_X1 rd_ptr_reg_25_ ( .D(n1521), .CLK(clk), .SN(1'b1), .Q(rd_ptr[25])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_26_ ( .D(n1581), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[26]) );
  DFFSNQ_X1 rd_ptr_reg_26_ ( .D(n1520), .CLK(clk), .SN(1'b1), .Q(rd_ptr[26])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_27_ ( .D(n1580), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[27]) );
  DFFSNQ_X1 rd_ptr_reg_27_ ( .D(n1519), .CLK(clk), .SN(1'b1), .Q(rd_ptr[27])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_28_ ( .D(n1579), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[28]) );
  DFFSNQ_X1 rd_ptr_reg_28_ ( .D(n1518), .CLK(clk), .SN(1'b1), .Q(rd_ptr[28])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_29_ ( .D(n1578), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[29]) );
  DFFSNQ_X1 rd_ptr_reg_29_ ( .D(n1517), .CLK(clk), .SN(1'b1), .Q(rd_ptr[29])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_30_ ( .D(n1577), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[30]) );
  DFFSNQ_X1 rd_ptr_reg_30_ ( .D(n1516), .CLK(clk), .SN(1'b1), .Q(rd_ptr[30])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_31_ ( .D(n1576), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[31]) );
  DFFSNQ_X1 rd_ptr_reg_31_ ( .D(n1515), .CLK(clk), .SN(1'b1), .Q(rd_ptr[31])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_32_ ( .D(n1575), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[32]) );
  DFFSNQ_X1 rd_ptr_reg_32_ ( .D(n1514), .CLK(clk), .SN(1'b1), .Q(rd_ptr[32])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_33_ ( .D(n1574), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[33]) );
  DFFSNQ_X1 rd_ptr_reg_33_ ( .D(n1513), .CLK(clk), .SN(1'b1), .Q(rd_ptr[33])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_34_ ( .D(n1573), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[34]) );
  DFFSNQ_X1 rd_ptr_reg_34_ ( .D(n1512), .CLK(clk), .SN(1'b1), .Q(rd_ptr[34])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_35_ ( .D(n1572), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[35]) );
  DFFSNQ_X1 rd_ptr_reg_35_ ( .D(n1511), .CLK(clk), .SN(1'b1), .Q(rd_ptr[35])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_36_ ( .D(n1571), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[36]) );
  DFFSNQ_X1 rd_ptr_reg_36_ ( .D(n1510), .CLK(clk), .SN(1'b1), .Q(rd_ptr[36])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_37_ ( .D(n1570), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[37]) );
  DFFSNQ_X1 rd_ptr_reg_37_ ( .D(n1509), .CLK(clk), .SN(1'b1), .Q(rd_ptr[37])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_38_ ( .D(n1569), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[38]) );
  DFFSNQ_X1 rd_ptr_reg_38_ ( .D(n1508), .CLK(clk), .SN(1'b1), .Q(rd_ptr[38])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_39_ ( .D(n1568), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[39]) );
  DFFSNQ_X1 rd_ptr_reg_39_ ( .D(n1507), .CLK(clk), .SN(1'b1), .Q(rd_ptr[39])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_40_ ( .D(n1567), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[40]) );
  DFFSNQ_X1 rd_ptr_reg_40_ ( .D(n1506), .CLK(clk), .SN(1'b1), .Q(rd_ptr[40])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_41_ ( .D(n1566), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[41]) );
  DFFSNQ_X1 rd_ptr_reg_41_ ( .D(n1505), .CLK(clk), .SN(1'b1), .Q(rd_ptr[41])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_42_ ( .D(n1565), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[42]) );
  DFFSNQ_X1 rd_ptr_reg_42_ ( .D(n1504), .CLK(clk), .SN(1'b1), .Q(rd_ptr[42])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_43_ ( .D(n1564), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[43]) );
  DFFSNQ_X1 rd_ptr_reg_43_ ( .D(n1503), .CLK(clk), .SN(1'b1), .Q(rd_ptr[43])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_44_ ( .D(n1563), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[44]) );
  DFFSNQ_X1 rd_ptr_reg_44_ ( .D(n1502), .CLK(clk), .SN(1'b1), .Q(rd_ptr[44])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_45_ ( .D(n1562), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[45]) );
  DFFSNQ_X1 rd_ptr_reg_45_ ( .D(n1501), .CLK(clk), .SN(1'b1), .Q(rd_ptr[45])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_46_ ( .D(n1561), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[46]) );
  DFFSNQ_X1 rd_ptr_reg_46_ ( .D(n1500), .CLK(clk), .SN(1'b1), .Q(rd_ptr[46])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_47_ ( .D(n1560), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[47]) );
  DFFSNQ_X1 rd_ptr_reg_47_ ( .D(n1499), .CLK(clk), .SN(1'b1), .Q(rd_ptr[47])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_48_ ( .D(n1559), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[48]) );
  DFFSNQ_X1 rd_ptr_reg_48_ ( .D(n1498), .CLK(clk), .SN(1'b1), .Q(rd_ptr[48])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_49_ ( .D(n1558), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[49]) );
  DFFSNQ_X1 rd_ptr_reg_49_ ( .D(n1497), .CLK(clk), .SN(1'b1), .Q(rd_ptr[49])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_50_ ( .D(n1557), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[50]) );
  DFFSNQ_X1 rd_ptr_reg_50_ ( .D(n1496), .CLK(clk), .SN(1'b1), .Q(rd_ptr[50])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_51_ ( .D(n1556), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[51]) );
  DFFSNQ_X1 rd_ptr_reg_51_ ( .D(n1495), .CLK(clk), .SN(1'b1), .Q(rd_ptr[51])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_52_ ( .D(n1555), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[52]) );
  DFFSNQ_X1 rd_ptr_reg_52_ ( .D(n1494), .CLK(clk), .SN(1'b1), .Q(rd_ptr[52])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_53_ ( .D(n1554), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[53]) );
  DFFSNQ_X1 rd_ptr_reg_53_ ( .D(n1493), .CLK(clk), .SN(1'b1), .Q(rd_ptr[53])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_54_ ( .D(n1553), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[54]) );
  DFFSNQ_X1 rd_ptr_reg_54_ ( .D(n1492), .CLK(clk), .SN(1'b1), .Q(rd_ptr[54])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_55_ ( .D(n1552), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[55]) );
  DFFSNQ_X1 rd_ptr_reg_55_ ( .D(n1491), .CLK(clk), .SN(1'b1), .Q(rd_ptr[55])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_56_ ( .D(n1551), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[56]) );
  DFFSNQ_X1 rd_ptr_reg_56_ ( .D(n1490), .CLK(clk), .SN(1'b1), .Q(rd_ptr[56])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_57_ ( .D(n1550), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[57]) );
  DFFSNQ_X1 rd_ptr_reg_57_ ( .D(n1489), .CLK(clk), .SN(1'b1), .Q(rd_ptr[57])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_58_ ( .D(n1549), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[58]) );
  DFFSNQ_X1 rd_ptr_reg_58_ ( .D(n1488), .CLK(clk), .SN(1'b1), .Q(rd_ptr[58])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_59_ ( .D(n1548), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[59]) );
  DFFSNQ_X1 rd_ptr_reg_59_ ( .D(n1487), .CLK(clk), .SN(1'b1), .Q(rd_ptr[59])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_60_ ( .D(n1547), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[60]) );
  DFFSNQ_X1 rd_ptr_reg_60_ ( .D(n1486), .CLK(clk), .SN(1'b1), .Q(rd_ptr[60])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_61_ ( .D(n1546), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[61]) );
  DFFSNQ_X1 rd_ptr_reg_61_ ( .D(n1485), .CLK(clk), .SN(1'b1), .Q(rd_ptr[61])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_62_ ( .D(n1545), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[62]) );
  DFFSNQ_X1 rd_ptr_reg_62_ ( .D(n1484), .CLK(clk), .SN(1'b1), .Q(rd_ptr[62])
         );
  DFFSNQ_X1 rd_ptr_reg_63_ ( .D(n1483), .CLK(clk), .SN(1'b1), .Q(rd_ptr[63])
         );
  DFFSNQ_X1 full_reg ( .D(n1482), .CLK(clk), .SN(1'b1), .Q(full) );
  DFFSNQ_X1 wr_ptr_reg_0_ ( .D(n1481), .CLK(clk), .SN(1'b1), .Q(wr_ptr[0]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_1_ ( .D(n642), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[1]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_2_ ( .D(n641), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[2]) );
  DFFSNQ_X1 wr_ptr_reg_2_ ( .D(n948), .CLK(clk), .SN(1'b1), .Q(wr_ptr[2]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_3_ ( .D(n640), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[3]) );
  DFFSNQ_X1 wr_ptr_reg_3_ ( .D(n947), .CLK(clk), .SN(1'b1), .Q(wr_ptr[3]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_4_ ( .D(n639), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[4]) );
  DFFSNQ_X1 wr_ptr_reg_4_ ( .D(n1480), .CLK(clk), .SN(1'b1), .Q(wr_ptr[4]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_5_ ( .D(n638), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[5]) );
  DFFSNQ_X1 wr_ptr_reg_5_ ( .D(n946), .CLK(clk), .SN(1'b1), .Q(wr_ptr[5]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_6_ ( .D(n637), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[6]) );
  DFFSNQ_X1 wr_ptr_reg_6_ ( .D(n945), .CLK(clk), .SN(1'b1), .Q(wr_ptr[6]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_7_ ( .D(n636), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[7]) );
  DFFSNQ_X1 wr_ptr_reg_7_ ( .D(n944), .CLK(clk), .SN(1'b1), .Q(wr_ptr[7]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_8_ ( .D(n635), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[8]) );
  DFFSNQ_X1 wr_ptr_reg_8_ ( .D(n943), .CLK(clk), .SN(1'b1), .Q(wr_ptr[8]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_9_ ( .D(n634), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[9]) );
  DFFSNQ_X1 wr_ptr_reg_9_ ( .D(n942), .CLK(clk), .SN(1'b1), .Q(wr_ptr[9]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_10_ ( .D(n633), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[10]) );
  DFFSNQ_X1 wr_ptr_reg_10_ ( .D(n1479), .CLK(clk), .SN(1'b1), .Q(wr_ptr[10])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_11_ ( .D(n632), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[11]) );
  DFFSNQ_X1 wr_ptr_reg_11_ ( .D(n1478), .CLK(clk), .SN(1'b1), .Q(wr_ptr[11])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_12_ ( .D(n631), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[12]) );
  DFFSNQ_X1 wr_ptr_reg_12_ ( .D(n1477), .CLK(clk), .SN(1'b1), .Q(wr_ptr[12])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_13_ ( .D(n630), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[13]) );
  DFFSNQ_X1 wr_ptr_reg_13_ ( .D(n941), .CLK(clk), .SN(1'b1), .Q(wr_ptr[13]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_14_ ( .D(n629), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[14]) );
  DFFSNQ_X1 wr_ptr_reg_14_ ( .D(n940), .CLK(clk), .SN(1'b1), .Q(wr_ptr[14]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_15_ ( .D(n628), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[15]) );
  DFFSNQ_X1 wr_ptr_reg_15_ ( .D(n939), .CLK(clk), .SN(1'b1), .Q(wr_ptr[15]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_16_ ( .D(n627), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[16]) );
  DFFSNQ_X1 wr_ptr_reg_16_ ( .D(n938), .CLK(clk), .SN(1'b1), .Q(wr_ptr[16]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_17_ ( .D(n626), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[17]) );
  DFFSNQ_X1 wr_ptr_reg_17_ ( .D(n937), .CLK(clk), .SN(1'b1), .Q(wr_ptr[17]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_18_ ( .D(n625), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[18]) );
  DFFSNQ_X1 wr_ptr_reg_18_ ( .D(n936), .CLK(clk), .SN(1'b1), .Q(wr_ptr[18]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_19_ ( .D(n624), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[19]) );
  DFFSNQ_X1 wr_ptr_reg_19_ ( .D(n935), .CLK(clk), .SN(1'b1), .Q(wr_ptr[19]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_20_ ( .D(n623), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[20]) );
  DFFSNQ_X1 wr_ptr_reg_20_ ( .D(n934), .CLK(clk), .SN(1'b1), .Q(wr_ptr[20]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_21_ ( .D(n622), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[21]) );
  DFFSNQ_X1 wr_ptr_reg_21_ ( .D(n933), .CLK(clk), .SN(1'b1), .Q(wr_ptr[21]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_22_ ( .D(n621), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[22]) );
  DFFSNQ_X1 wr_ptr_reg_22_ ( .D(n932), .CLK(clk), .SN(1'b1), .Q(wr_ptr[22]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_23_ ( .D(n620), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[23]) );
  DFFSNQ_X1 wr_ptr_reg_23_ ( .D(n931), .CLK(clk), .SN(1'b1), .Q(wr_ptr[23]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_24_ ( .D(n619), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[24]) );
  DFFSNQ_X1 wr_ptr_reg_24_ ( .D(n930), .CLK(clk), .SN(1'b1), .Q(wr_ptr[24]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_25_ ( .D(n618), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[25]) );
  DFFSNQ_X1 wr_ptr_reg_25_ ( .D(n929), .CLK(clk), .SN(1'b1), .Q(wr_ptr[25]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_26_ ( .D(n617), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[26]) );
  DFFSNQ_X1 wr_ptr_reg_26_ ( .D(n928), .CLK(clk), .SN(1'b1), .Q(wr_ptr[26]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_27_ ( .D(n616), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[27]) );
  DFFSNQ_X1 wr_ptr_reg_27_ ( .D(n927), .CLK(clk), .SN(1'b1), .Q(wr_ptr[27]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_28_ ( .D(n615), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[28]) );
  DFFSNQ_X1 wr_ptr_reg_28_ ( .D(n926), .CLK(clk), .SN(1'b1), .Q(wr_ptr[28]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_29_ ( .D(n614), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[29]) );
  DFFSNQ_X1 wr_ptr_reg_29_ ( .D(n925), .CLK(clk), .SN(1'b1), .Q(wr_ptr[29]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_30_ ( .D(n613), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[30]) );
  DFFSNQ_X1 wr_ptr_reg_30_ ( .D(n924), .CLK(clk), .SN(1'b1), .Q(wr_ptr[30]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_31_ ( .D(n612), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[31]) );
  DFFSNQ_X1 wr_ptr_reg_31_ ( .D(n923), .CLK(clk), .SN(1'b1), .Q(wr_ptr[31]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_32_ ( .D(n611), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[32]) );
  DFFSNQ_X1 wr_ptr_reg_32_ ( .D(n922), .CLK(clk), .SN(1'b1), .Q(wr_ptr[32]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_33_ ( .D(n610), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[33]) );
  DFFSNQ_X1 wr_ptr_reg_33_ ( .D(n921), .CLK(clk), .SN(1'b1), .Q(wr_ptr[33]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_34_ ( .D(n609), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[34]) );
  DFFSNQ_X1 wr_ptr_reg_34_ ( .D(n920), .CLK(clk), .SN(1'b1), .Q(wr_ptr[34]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_35_ ( .D(n608), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[35]) );
  DFFSNQ_X1 wr_ptr_reg_35_ ( .D(n919), .CLK(clk), .SN(1'b1), .Q(wr_ptr[35]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_36_ ( .D(n607), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[36]) );
  DFFSNQ_X1 wr_ptr_reg_36_ ( .D(n918), .CLK(clk), .SN(1'b1), .Q(wr_ptr[36]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_37_ ( .D(n606), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[37]) );
  DFFSNQ_X1 wr_ptr_reg_37_ ( .D(n917), .CLK(clk), .SN(1'b1), .Q(wr_ptr[37]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_38_ ( .D(n605), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[38]) );
  DFFSNQ_X1 wr_ptr_reg_38_ ( .D(n916), .CLK(clk), .SN(1'b1), .Q(wr_ptr[38]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_39_ ( .D(n604), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[39]) );
  DFFSNQ_X1 wr_ptr_reg_39_ ( .D(n915), .CLK(clk), .SN(1'b1), .Q(wr_ptr[39]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_40_ ( .D(n603), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[40]) );
  DFFSNQ_X1 wr_ptr_reg_40_ ( .D(n914), .CLK(clk), .SN(1'b1), .Q(wr_ptr[40]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_41_ ( .D(n602), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[41]) );
  DFFSNQ_X1 wr_ptr_reg_41_ ( .D(n913), .CLK(clk), .SN(1'b1), .Q(wr_ptr[41]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_42_ ( .D(n601), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[42]) );
  DFFSNQ_X1 wr_ptr_reg_42_ ( .D(n912), .CLK(clk), .SN(1'b1), .Q(wr_ptr[42]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_43_ ( .D(n600), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[43]) );
  DFFSNQ_X1 wr_ptr_reg_43_ ( .D(n911), .CLK(clk), .SN(1'b1), .Q(wr_ptr[43]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_44_ ( .D(n599), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[44]) );
  DFFSNQ_X1 wr_ptr_reg_44_ ( .D(n910), .CLK(clk), .SN(1'b1), .Q(wr_ptr[44]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_45_ ( .D(n598), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[45]) );
  DFFSNQ_X1 wr_ptr_reg_45_ ( .D(n909), .CLK(clk), .SN(1'b1), .Q(wr_ptr[45]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_46_ ( .D(n597), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[46]) );
  DFFSNQ_X1 wr_ptr_reg_46_ ( .D(n1476), .CLK(clk), .SN(1'b1), .Q(wr_ptr[46])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_47_ ( .D(n596), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[47]) );
  DFFSNQ_X1 wr_ptr_reg_47_ ( .D(n1475), .CLK(clk), .SN(1'b1), .Q(wr_ptr[47])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_48_ ( .D(n595), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[48]) );
  DFFSNQ_X1 wr_ptr_reg_48_ ( .D(n1474), .CLK(clk), .SN(1'b1), .Q(wr_ptr[48])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_49_ ( .D(n594), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[49]) );
  DFFSNQ_X1 wr_ptr_reg_49_ ( .D(n1473), .CLK(clk), .SN(1'b1), .Q(wr_ptr[49])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_50_ ( .D(n593), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[50]) );
  DFFSNQ_X1 wr_ptr_reg_50_ ( .D(n1472), .CLK(clk), .SN(1'b1), .Q(wr_ptr[50])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_51_ ( .D(n592), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[51]) );
  DFFSNQ_X1 wr_ptr_reg_51_ ( .D(n1471), .CLK(clk), .SN(1'b1), .Q(wr_ptr[51])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_52_ ( .D(n591), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[52]) );
  DFFSNQ_X1 wr_ptr_reg_52_ ( .D(n1470), .CLK(clk), .SN(1'b1), .Q(wr_ptr[52])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_53_ ( .D(n590), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[53]) );
  DFFSNQ_X1 wr_ptr_reg_53_ ( .D(n908), .CLK(clk), .SN(1'b1), .Q(wr_ptr[53]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_54_ ( .D(n589), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[54]) );
  DFFSNQ_X1 wr_ptr_reg_54_ ( .D(n907), .CLK(clk), .SN(1'b1), .Q(wr_ptr[54]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_55_ ( .D(n588), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[55]) );
  DFFSNQ_X1 wr_ptr_reg_55_ ( .D(n906), .CLK(clk), .SN(1'b1), .Q(wr_ptr[55]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_56_ ( .D(n587), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[56]) );
  DFFSNQ_X1 wr_ptr_reg_56_ ( .D(n905), .CLK(clk), .SN(1'b1), .Q(wr_ptr[56]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_57_ ( .D(n586), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[57]) );
  DFFSNQ_X1 wr_ptr_reg_57_ ( .D(n904), .CLK(clk), .SN(1'b1), .Q(wr_ptr[57]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_58_ ( .D(n585), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[58]) );
  DFFSNQ_X1 wr_ptr_reg_58_ ( .D(n903), .CLK(clk), .SN(1'b1), .Q(wr_ptr[58]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_59_ ( .D(n584), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[59]) );
  DFFSNQ_X1 wr_ptr_reg_59_ ( .D(n902), .CLK(clk), .SN(1'b1), .Q(wr_ptr[59]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_60_ ( .D(n583), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[60]) );
  DFFSNQ_X1 wr_ptr_reg_60_ ( .D(n901), .CLK(clk), .SN(1'b1), .Q(wr_ptr[60]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_61_ ( .D(n582), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[61]) );
  DFFSNQ_X1 wr_ptr_reg_61_ ( .D(n900), .CLK(clk), .SN(1'b1), .Q(wr_ptr[61]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_62_ ( .D(n581), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[62]) );
  DFFSNQ_X1 wr_ptr_reg_62_ ( .D(n899), .CLK(clk), .SN(1'b1), .Q(wr_ptr[62]) );
  DFFSNQ_X1 wr_ptr_reg_1_ ( .D(n949), .CLK(clk), .SN(1'b1), .Q(wr_ptr[1]) );
  DFFSNQ_X1 wr_ptr_reg_63_ ( .D(n644), .CLK(clk), .SN(1'b1), .Q(wr_ptr[63]) );
  DFFSNQ_X1 queue_reg_1__63_ ( .D(n1648), .CLK(clk), .SN(1'b1), .Q(queue[127])
         );
  DFFSNQ_X1 queue_reg_1__62_ ( .D(n1649), .CLK(clk), .SN(1'b1), .Q(queue[126])
         );
  DFFSNQ_X1 queue_reg_1__61_ ( .D(n1650), .CLK(clk), .SN(1'b1), .Q(queue[125])
         );
  DFFSNQ_X1 queue_reg_1__60_ ( .D(n1651), .CLK(clk), .SN(1'b1), .Q(queue[124])
         );
  DFFSNQ_X1 queue_reg_1__59_ ( .D(n1652), .CLK(clk), .SN(1'b1), .Q(queue[123])
         );
  DFFSNQ_X1 queue_reg_1__58_ ( .D(n1653), .CLK(clk), .SN(1'b1), .Q(queue[122])
         );
  DFFSNQ_X1 queue_reg_1__57_ ( .D(n1654), .CLK(clk), .SN(1'b1), .Q(queue[121])
         );
  DFFSNQ_X1 queue_reg_1__56_ ( .D(n1655), .CLK(clk), .SN(1'b1), .Q(queue[120])
         );
  DFFSNQ_X1 queue_reg_1__55_ ( .D(n1656), .CLK(clk), .SN(1'b1), .Q(queue[119])
         );
  DFFSNQ_X1 queue_reg_1__54_ ( .D(n1657), .CLK(clk), .SN(1'b1), .Q(queue[118])
         );
  DFFSNQ_X1 queue_reg_1__53_ ( .D(n1658), .CLK(clk), .SN(1'b1), .Q(queue[117])
         );
  DFFSNQ_X1 queue_reg_1__52_ ( .D(n1659), .CLK(clk), .SN(1'b1), .Q(queue[116])
         );
  DFFSNQ_X1 queue_reg_1__51_ ( .D(n1660), .CLK(clk), .SN(1'b1), .Q(queue[115])
         );
  DFFSNQ_X1 queue_reg_1__50_ ( .D(n1661), .CLK(clk), .SN(1'b1), .Q(queue[114])
         );
  DFFSNQ_X1 queue_reg_1__49_ ( .D(n1662), .CLK(clk), .SN(1'b1), .Q(queue[113])
         );
  DFFSNQ_X1 queue_reg_1__48_ ( .D(n1663), .CLK(clk), .SN(1'b1), .Q(queue[112])
         );
  DFFSNQ_X1 queue_reg_1__47_ ( .D(n1664), .CLK(clk), .SN(1'b1), .Q(queue[111])
         );
  DFFSNQ_X1 queue_reg_1__46_ ( .D(n1665), .CLK(clk), .SN(1'b1), .Q(queue[110])
         );
  DFFSNQ_X1 queue_reg_1__45_ ( .D(n1666), .CLK(clk), .SN(1'b1), .Q(queue[109])
         );
  DFFSNQ_X1 queue_reg_1__44_ ( .D(n1667), .CLK(clk), .SN(1'b1), .Q(queue[108])
         );
  DFFSNQ_X1 queue_reg_1__43_ ( .D(n1668), .CLK(clk), .SN(1'b1), .Q(queue[107])
         );
  DFFSNQ_X1 queue_reg_1__42_ ( .D(n1669), .CLK(clk), .SN(1'b1), .Q(queue[106])
         );
  DFFSNQ_X1 queue_reg_1__41_ ( .D(n1670), .CLK(clk), .SN(1'b1), .Q(queue[105])
         );
  DFFSNQ_X1 queue_reg_1__40_ ( .D(n1671), .CLK(clk), .SN(1'b1), .Q(queue[104])
         );
  DFFSNQ_X1 queue_reg_1__39_ ( .D(n1672), .CLK(clk), .SN(1'b1), .Q(queue[103])
         );
  DFFSNQ_X1 queue_reg_1__38_ ( .D(n1673), .CLK(clk), .SN(1'b1), .Q(queue[102])
         );
  DFFSNQ_X1 queue_reg_1__37_ ( .D(n1674), .CLK(clk), .SN(1'b1), .Q(queue[101])
         );
  DFFSNQ_X1 queue_reg_1__36_ ( .D(n1675), .CLK(clk), .SN(1'b1), .Q(queue[100])
         );
  DFFSNQ_X1 queue_reg_1__35_ ( .D(n1676), .CLK(clk), .SN(1'b1), .Q(queue[99])
         );
  DFFSNQ_X1 queue_reg_1__34_ ( .D(n1677), .CLK(clk), .SN(1'b1), .Q(queue[98])
         );
  DFFSNQ_X1 queue_reg_1__33_ ( .D(n1678), .CLK(clk), .SN(1'b1), .Q(queue[97])
         );
  DFFSNQ_X1 queue_reg_1__32_ ( .D(n1679), .CLK(clk), .SN(1'b1), .Q(queue[96])
         );
  DFFSNQ_X1 queue_reg_1__31_ ( .D(n1680), .CLK(clk), .SN(1'b1), .Q(queue[95])
         );
  DFFSNQ_X1 queue_reg_1__30_ ( .D(n1681), .CLK(clk), .SN(1'b1), .Q(queue[94])
         );
  DFFSNQ_X1 queue_reg_1__29_ ( .D(n1682), .CLK(clk), .SN(1'b1), .Q(queue[93])
         );
  DFFSNQ_X1 queue_reg_1__28_ ( .D(n1683), .CLK(clk), .SN(1'b1), .Q(queue[92])
         );
  DFFSNQ_X1 queue_reg_1__27_ ( .D(n1684), .CLK(clk), .SN(1'b1), .Q(queue[91])
         );
  DFFSNQ_X1 queue_reg_1__26_ ( .D(n1685), .CLK(clk), .SN(1'b1), .Q(queue[90])
         );
  DFFSNQ_X1 queue_reg_1__25_ ( .D(n1686), .CLK(clk), .SN(1'b1), .Q(queue[89])
         );
  DFFSNQ_X1 queue_reg_1__24_ ( .D(n1687), .CLK(clk), .SN(1'b1), .Q(queue[88])
         );
  DFFSNQ_X1 queue_reg_1__23_ ( .D(n1688), .CLK(clk), .SN(1'b1), .Q(queue[87])
         );
  DFFSNQ_X1 queue_reg_1__22_ ( .D(n1689), .CLK(clk), .SN(1'b1), .Q(queue[86])
         );
  DFFSNQ_X1 queue_reg_1__21_ ( .D(n1690), .CLK(clk), .SN(1'b1), .Q(queue[85])
         );
  DFFSNQ_X1 queue_reg_1__20_ ( .D(n1691), .CLK(clk), .SN(1'b1), .Q(queue[84])
         );
  DFFSNQ_X1 queue_reg_1__19_ ( .D(n1692), .CLK(clk), .SN(1'b1), .Q(queue[83])
         );
  DFFSNQ_X1 queue_reg_1__18_ ( .D(n1693), .CLK(clk), .SN(1'b1), .Q(queue[82])
         );
  DFFSNQ_X1 queue_reg_1__17_ ( .D(n1694), .CLK(clk), .SN(1'b1), .Q(queue[81])
         );
  DFFSNQ_X1 queue_reg_1__16_ ( .D(n1695), .CLK(clk), .SN(1'b1), .Q(queue[80])
         );
  DFFSNQ_X1 queue_reg_1__15_ ( .D(n1696), .CLK(clk), .SN(1'b1), .Q(queue[79])
         );
  DFFSNQ_X1 queue_reg_1__14_ ( .D(n1697), .CLK(clk), .SN(1'b1), .Q(queue[78])
         );
  DFFSNQ_X1 queue_reg_1__13_ ( .D(n1698), .CLK(clk), .SN(1'b1), .Q(queue[77])
         );
  DFFSNQ_X1 queue_reg_1__12_ ( .D(n1699), .CLK(clk), .SN(1'b1), .Q(queue[76])
         );
  DFFSNQ_X1 queue_reg_1__11_ ( .D(n1700), .CLK(clk), .SN(1'b1), .Q(queue[75])
         );
  DFFSNQ_X1 queue_reg_1__10_ ( .D(n1701), .CLK(clk), .SN(1'b1), .Q(queue[74])
         );
  DFFSNQ_X1 queue_reg_1__9_ ( .D(n1702), .CLK(clk), .SN(1'b1), .Q(queue[73])
         );
  DFFSNQ_X1 queue_reg_1__8_ ( .D(n1703), .CLK(clk), .SN(1'b1), .Q(queue[72])
         );
  DFFSNQ_X1 queue_reg_1__7_ ( .D(n1704), .CLK(clk), .SN(1'b1), .Q(queue[71])
         );
  DFFSNQ_X1 queue_reg_1__6_ ( .D(n1705), .CLK(clk), .SN(1'b1), .Q(queue[70])
         );
  DFFSNQ_X1 queue_reg_1__5_ ( .D(n1706), .CLK(clk), .SN(1'b1), .Q(queue[69])
         );
  DFFSNQ_X1 queue_reg_1__4_ ( .D(n1707), .CLK(clk), .SN(1'b1), .Q(queue[68])
         );
  DFFSNQ_X1 queue_reg_1__3_ ( .D(n1708), .CLK(clk), .SN(1'b1), .Q(queue[67])
         );
  DFFSNQ_X1 queue_reg_1__2_ ( .D(n1709), .CLK(clk), .SN(1'b1), .Q(queue[66])
         );
  DFFSNQ_X1 queue_reg_1__1_ ( .D(n1710), .CLK(clk), .SN(1'b1), .Q(queue[65])
         );
  DFFSNQ_X1 queue_reg_1__0_ ( .D(n1711), .CLK(clk), .SN(1'b1), .Q(queue[64])
         );
  DFFSNQ_X1 queue_reg_0__63_ ( .D(n951), .CLK(clk), .SN(1'b1), .Q(queue[63])
         );
  DFFSNQ_X1 queue_reg_0__62_ ( .D(n952), .CLK(clk), .SN(1'b1), .Q(queue[62])
         );
  DFFSNQ_X1 queue_reg_0__61_ ( .D(n953), .CLK(clk), .SN(1'b1), .Q(queue[61])
         );
  DFFSNQ_X1 queue_reg_0__60_ ( .D(n954), .CLK(clk), .SN(1'b1), .Q(queue[60])
         );
  DFFSNQ_X1 queue_reg_0__59_ ( .D(n955), .CLK(clk), .SN(1'b1), .Q(queue[59])
         );
  DFFSNQ_X1 queue_reg_0__58_ ( .D(n956), .CLK(clk), .SN(1'b1), .Q(queue[58])
         );
  DFFSNQ_X1 queue_reg_0__57_ ( .D(n957), .CLK(clk), .SN(1'b1), .Q(queue[57])
         );
  DFFSNQ_X1 queue_reg_0__56_ ( .D(n958), .CLK(clk), .SN(1'b1), .Q(queue[56])
         );
  DFFSNQ_X1 queue_reg_0__55_ ( .D(n959), .CLK(clk), .SN(1'b1), .Q(queue[55])
         );
  DFFSNQ_X1 queue_reg_0__54_ ( .D(n960), .CLK(clk), .SN(1'b1), .Q(queue[54])
         );
  DFFSNQ_X1 queue_reg_0__53_ ( .D(n961), .CLK(clk), .SN(1'b1), .Q(queue[53])
         );
  DFFSNQ_X1 queue_reg_0__52_ ( .D(n962), .CLK(clk), .SN(1'b1), .Q(queue[52])
         );
  DFFSNQ_X1 queue_reg_0__51_ ( .D(n963), .CLK(clk), .SN(1'b1), .Q(queue[51])
         );
  DFFSNQ_X1 queue_reg_0__50_ ( .D(n964), .CLK(clk), .SN(1'b1), .Q(queue[50])
         );
  DFFSNQ_X1 queue_reg_0__49_ ( .D(n965), .CLK(clk), .SN(1'b1), .Q(queue[49])
         );
  DFFSNQ_X1 queue_reg_0__48_ ( .D(n966), .CLK(clk), .SN(1'b1), .Q(queue[48])
         );
  DFFSNQ_X1 queue_reg_0__47_ ( .D(n967), .CLK(clk), .SN(1'b1), .Q(queue[47])
         );
  DFFSNQ_X1 queue_reg_0__46_ ( .D(n968), .CLK(clk), .SN(1'b1), .Q(queue[46])
         );
  DFFSNQ_X1 queue_reg_0__45_ ( .D(n969), .CLK(clk), .SN(1'b1), .Q(queue[45])
         );
  DFFSNQ_X1 queue_reg_0__44_ ( .D(n970), .CLK(clk), .SN(1'b1), .Q(queue[44])
         );
  DFFSNQ_X1 queue_reg_0__43_ ( .D(n971), .CLK(clk), .SN(1'b1), .Q(queue[43])
         );
  DFFSNQ_X1 queue_reg_0__42_ ( .D(n972), .CLK(clk), .SN(1'b1), .Q(queue[42])
         );
  DFFSNQ_X1 queue_reg_0__41_ ( .D(n973), .CLK(clk), .SN(1'b1), .Q(queue[41])
         );
  DFFSNQ_X1 queue_reg_0__40_ ( .D(n974), .CLK(clk), .SN(1'b1), .Q(queue[40])
         );
  DFFSNQ_X1 queue_reg_0__39_ ( .D(n975), .CLK(clk), .SN(1'b1), .Q(queue[39])
         );
  DFFSNQ_X1 queue_reg_0__38_ ( .D(n976), .CLK(clk), .SN(1'b1), .Q(queue[38])
         );
  DFFSNQ_X1 queue_reg_0__37_ ( .D(n1336), .CLK(clk), .SN(1'b1), .Q(queue[37])
         );
  DFFSNQ_X1 queue_reg_0__36_ ( .D(n1611), .CLK(clk), .SN(1'b1), .Q(queue[36])
         );
  DFFSNQ_X1 queue_reg_0__35_ ( .D(n1612), .CLK(clk), .SN(1'b1), .Q(queue[35])
         );
  DFFSNQ_X1 queue_reg_0__34_ ( .D(n1613), .CLK(clk), .SN(1'b1), .Q(queue[34])
         );
  DFFSNQ_X1 queue_reg_0__33_ ( .D(n1614), .CLK(clk), .SN(1'b1), .Q(queue[33])
         );
  DFFSNQ_X1 queue_reg_0__32_ ( .D(n1615), .CLK(clk), .SN(1'b1), .Q(queue[32])
         );
  DFFSNQ_X1 queue_reg_0__31_ ( .D(n1616), .CLK(clk), .SN(1'b1), .Q(queue[31])
         );
  DFFSNQ_X1 queue_reg_0__30_ ( .D(n1617), .CLK(clk), .SN(1'b1), .Q(queue[30])
         );
  DFFSNQ_X1 queue_reg_0__29_ ( .D(n1618), .CLK(clk), .SN(1'b1), .Q(queue[29])
         );
  DFFSNQ_X1 queue_reg_0__28_ ( .D(n1619), .CLK(clk), .SN(1'b1), .Q(queue[28])
         );
  DFFSNQ_X1 queue_reg_0__27_ ( .D(n1620), .CLK(clk), .SN(1'b1), .Q(queue[27])
         );
  DFFSNQ_X1 queue_reg_0__26_ ( .D(n1621), .CLK(clk), .SN(1'b1), .Q(queue[26])
         );
  DFFSNQ_X1 queue_reg_0__25_ ( .D(n1622), .CLK(clk), .SN(1'b1), .Q(queue[25])
         );
  DFFSNQ_X1 queue_reg_0__24_ ( .D(n1623), .CLK(clk), .SN(1'b1), .Q(queue[24])
         );
  DFFSNQ_X1 queue_reg_0__23_ ( .D(n1624), .CLK(clk), .SN(1'b1), .Q(queue[23])
         );
  DFFSNQ_X1 queue_reg_0__22_ ( .D(n1625), .CLK(clk), .SN(1'b1), .Q(queue[22])
         );
  DFFSNQ_X1 queue_reg_0__21_ ( .D(n1626), .CLK(clk), .SN(1'b1), .Q(queue[21])
         );
  DFFSNQ_X1 queue_reg_0__20_ ( .D(n1627), .CLK(clk), .SN(1'b1), .Q(queue[20])
         );
  DFFSNQ_X1 queue_reg_0__19_ ( .D(n1628), .CLK(clk), .SN(1'b1), .Q(queue[19])
         );
  DFFSNQ_X1 queue_reg_0__18_ ( .D(n1629), .CLK(clk), .SN(1'b1), .Q(queue[18])
         );
  DFFSNQ_X1 queue_reg_0__17_ ( .D(n1630), .CLK(clk), .SN(1'b1), .Q(queue[17])
         );
  DFFSNQ_X1 queue_reg_0__16_ ( .D(n1631), .CLK(clk), .SN(1'b1), .Q(queue[16])
         );
  DFFSNQ_X1 queue_reg_0__15_ ( .D(n1632), .CLK(clk), .SN(1'b1), .Q(queue[15])
         );
  DFFSNQ_X1 queue_reg_0__14_ ( .D(n1633), .CLK(clk), .SN(1'b1), .Q(queue[14])
         );
  DFFSNQ_X1 queue_reg_0__13_ ( .D(n1634), .CLK(clk), .SN(1'b1), .Q(queue[13])
         );
  DFFSNQ_X1 queue_reg_0__12_ ( .D(n1635), .CLK(clk), .SN(1'b1), .Q(queue[12])
         );
  DFFSNQ_X1 queue_reg_0__11_ ( .D(n1636), .CLK(clk), .SN(1'b1), .Q(queue[11])
         );
  DFFSNQ_X1 queue_reg_0__10_ ( .D(n1637), .CLK(clk), .SN(1'b1), .Q(queue[10])
         );
  DFFSNQ_X1 queue_reg_0__9_ ( .D(n1638), .CLK(clk), .SN(1'b1), .Q(queue[9]) );
  DFFSNQ_X1 queue_reg_0__8_ ( .D(n1639), .CLK(clk), .SN(1'b1), .Q(queue[8]) );
  DFFSNQ_X1 queue_reg_0__7_ ( .D(n1640), .CLK(clk), .SN(1'b1), .Q(queue[7]) );
  DFFSNQ_X1 queue_reg_0__6_ ( .D(n1641), .CLK(clk), .SN(1'b1), .Q(queue[6]) );
  DFFSNQ_X1 queue_reg_0__5_ ( .D(n1642), .CLK(clk), .SN(1'b1), .Q(queue[5]) );
  DFFSNQ_X1 queue_reg_0__4_ ( .D(n1643), .CLK(clk), .SN(1'b1), .Q(queue[4]) );
  DFFSNQ_X1 queue_reg_0__3_ ( .D(n1644), .CLK(clk), .SN(1'b1), .Q(queue[3]) );
  DFFSNQ_X1 queue_reg_0__2_ ( .D(n1645), .CLK(clk), .SN(1'b1), .Q(queue[2]) );
  DFFSNQ_X1 queue_reg_0__1_ ( .D(n1646), .CLK(clk), .SN(1'b1), .Q(queue[1]) );
  DFFSNQ_X1 queue_reg_0__0_ ( .D(n1647), .CLK(clk), .SN(1'b1), .Q(queue[0]) );
  DFFSNQ_X1 data_out_reg_63_ ( .D(n645), .CLK(clk), .SN(1'b1), .Q(data_out[63]) );
  DFFSNQ_X1 data_out_reg_62_ ( .D(n646), .CLK(clk), .SN(1'b1), .Q(data_out[62]) );
  DFFSNQ_X1 data_out_reg_61_ ( .D(n647), .CLK(clk), .SN(1'b1), .Q(data_out[61]) );
  DFFSNQ_X1 data_out_reg_60_ ( .D(n648), .CLK(clk), .SN(1'b1), .Q(data_out[60]) );
  DFFSNQ_X1 data_out_reg_59_ ( .D(n649), .CLK(clk), .SN(1'b1), .Q(data_out[59]) );
  DFFSNQ_X1 data_out_reg_58_ ( .D(n650), .CLK(clk), .SN(1'b1), .Q(data_out[58]) );
  DFFSNQ_X1 data_out_reg_57_ ( .D(n651), .CLK(clk), .SN(1'b1), .Q(data_out[57]) );
  DFFSNQ_X1 data_out_reg_56_ ( .D(n652), .CLK(clk), .SN(1'b1), .Q(data_out[56]) );
  DFFSNQ_X1 data_out_reg_55_ ( .D(n653), .CLK(clk), .SN(1'b1), .Q(data_out[55]) );
  DFFSNQ_X1 data_out_reg_54_ ( .D(n654), .CLK(clk), .SN(1'b1), .Q(data_out[54]) );
  DFFSNQ_X1 data_out_reg_53_ ( .D(n655), .CLK(clk), .SN(1'b1), .Q(data_out[53]) );
  DFFSNQ_X1 data_out_reg_52_ ( .D(n656), .CLK(clk), .SN(1'b1), .Q(data_out[52]) );
  DFFSNQ_X1 data_out_reg_51_ ( .D(n657), .CLK(clk), .SN(1'b1), .Q(data_out[51]) );
  DFFSNQ_X1 data_out_reg_50_ ( .D(n658), .CLK(clk), .SN(1'b1), .Q(data_out[50]) );
  DFFSNQ_X1 data_out_reg_49_ ( .D(n659), .CLK(clk), .SN(1'b1), .Q(data_out[49]) );
  DFFSNQ_X1 data_out_reg_48_ ( .D(n660), .CLK(clk), .SN(1'b1), .Q(data_out[48]) );
  DFFSNQ_X1 data_out_reg_47_ ( .D(n661), .CLK(clk), .SN(1'b1), .Q(data_out[47]) );
  DFFSNQ_X1 data_out_reg_46_ ( .D(n662), .CLK(clk), .SN(1'b1), .Q(data_out[46]) );
  DFFSNQ_X1 data_out_reg_45_ ( .D(n663), .CLK(clk), .SN(1'b1), .Q(data_out[45]) );
  DFFSNQ_X1 data_out_reg_44_ ( .D(n664), .CLK(clk), .SN(1'b1), .Q(data_out[44]) );
  DFFSNQ_X1 data_out_reg_43_ ( .D(n665), .CLK(clk), .SN(1'b1), .Q(data_out[43]) );
  DFFSNQ_X1 data_out_reg_42_ ( .D(n666), .CLK(clk), .SN(1'b1), .Q(data_out[42]) );
  DFFSNQ_X1 data_out_reg_41_ ( .D(n667), .CLK(clk), .SN(1'b1), .Q(data_out[41]) );
  DFFSNQ_X1 data_out_reg_40_ ( .D(n668), .CLK(clk), .SN(1'b1), .Q(data_out[40]) );
  DFFSNQ_X1 data_out_reg_39_ ( .D(n669), .CLK(clk), .SN(1'b1), .Q(data_out[39]) );
  DFFSNQ_X1 data_out_reg_38_ ( .D(n670), .CLK(clk), .SN(1'b1), .Q(data_out[38]) );
  DFFSNQ_X1 data_out_reg_37_ ( .D(n671), .CLK(clk), .SN(1'b1), .Q(data_out[37]) );
  DFFSNQ_X1 data_out_reg_36_ ( .D(n672), .CLK(clk), .SN(1'b1), .Q(data_out[36]) );
  DFFSNQ_X1 data_out_reg_35_ ( .D(n673), .CLK(clk), .SN(1'b1), .Q(data_out[35]) );
  DFFSNQ_X1 data_out_reg_34_ ( .D(n674), .CLK(clk), .SN(1'b1), .Q(data_out[34]) );
  DFFSNQ_X1 data_out_reg_33_ ( .D(n675), .CLK(clk), .SN(1'b1), .Q(data_out[33]) );
  DFFSNQ_X1 data_out_reg_32_ ( .D(n676), .CLK(clk), .SN(1'b1), .Q(data_out[32]) );
  DFFSNQ_X1 data_out_reg_31_ ( .D(n677), .CLK(clk), .SN(1'b1), .Q(data_out[31]) );
  DFFSNQ_X1 data_out_reg_30_ ( .D(n678), .CLK(clk), .SN(1'b1), .Q(data_out[30]) );
  DFFSNQ_X1 data_out_reg_29_ ( .D(n679), .CLK(clk), .SN(1'b1), .Q(data_out[29]) );
  DFFSNQ_X1 data_out_reg_28_ ( .D(n680), .CLK(clk), .SN(1'b1), .Q(data_out[28]) );
  DFFSNQ_X1 data_out_reg_27_ ( .D(n681), .CLK(clk), .SN(1'b1), .Q(data_out[27]) );
  DFFSNQ_X1 data_out_reg_26_ ( .D(n682), .CLK(clk), .SN(1'b1), .Q(data_out[26]) );
  DFFSNQ_X1 data_out_reg_25_ ( .D(n683), .CLK(clk), .SN(1'b1), .Q(data_out[25]) );
  DFFSNQ_X1 data_out_reg_24_ ( .D(n684), .CLK(clk), .SN(1'b1), .Q(data_out[24]) );
  DFFSNQ_X1 data_out_reg_23_ ( .D(n685), .CLK(clk), .SN(1'b1), .Q(data_out[23]) );
  DFFSNQ_X1 data_out_reg_22_ ( .D(n686), .CLK(clk), .SN(1'b1), .Q(data_out[22]) );
  DFFSNQ_X1 data_out_reg_21_ ( .D(n687), .CLK(clk), .SN(1'b1), .Q(data_out[21]) );
  DFFSNQ_X1 data_out_reg_20_ ( .D(n688), .CLK(clk), .SN(1'b1), .Q(data_out[20]) );
  DFFSNQ_X1 data_out_reg_19_ ( .D(n689), .CLK(clk), .SN(1'b1), .Q(data_out[19]) );
  DFFSNQ_X1 data_out_reg_18_ ( .D(n690), .CLK(clk), .SN(1'b1), .Q(data_out[18]) );
  DFFSNQ_X1 data_out_reg_17_ ( .D(n691), .CLK(clk), .SN(1'b1), .Q(data_out[17]) );
  DFFSNQ_X1 data_out_reg_16_ ( .D(n692), .CLK(clk), .SN(1'b1), .Q(data_out[16]) );
  DFFSNQ_X1 data_out_reg_15_ ( .D(n693), .CLK(clk), .SN(1'b1), .Q(data_out[15]) );
  DFFSNQ_X1 data_out_reg_14_ ( .D(n694), .CLK(clk), .SN(1'b1), .Q(data_out[14]) );
  DFFSNQ_X1 data_out_reg_13_ ( .D(n695), .CLK(clk), .SN(1'b1), .Q(data_out[13]) );
  DFFSNQ_X1 data_out_reg_12_ ( .D(n696), .CLK(clk), .SN(1'b1), .Q(data_out[12]) );
  DFFSNQ_X1 data_out_reg_11_ ( .D(n697), .CLK(clk), .SN(1'b1), .Q(data_out[11]) );
  DFFSNQ_X1 data_out_reg_10_ ( .D(n698), .CLK(clk), .SN(1'b1), .Q(data_out[10]) );
  DFFSNQ_X1 data_out_reg_9_ ( .D(n699), .CLK(clk), .SN(1'b1), .Q(data_out[9])
         );
  DFFSNQ_X1 data_out_reg_8_ ( .D(n700), .CLK(clk), .SN(1'b1), .Q(data_out[8])
         );
  DFFSNQ_X1 data_out_reg_7_ ( .D(n701), .CLK(clk), .SN(1'b1), .Q(data_out[7])
         );
  DFFSNQ_X1 data_out_reg_6_ ( .D(n702), .CLK(clk), .SN(1'b1), .Q(data_out[6])
         );
  DFFSNQ_X1 data_out_reg_5_ ( .D(n703), .CLK(clk), .SN(1'b1), .Q(data_out[5])
         );
  DFFSNQ_X1 data_out_reg_4_ ( .D(n704), .CLK(clk), .SN(1'b1), .Q(data_out[4])
         );
  DFFSNQ_X1 data_out_reg_3_ ( .D(n705), .CLK(clk), .SN(1'b1), .Q(data_out[3])
         );
  DFFSNQ_X1 data_out_reg_2_ ( .D(n706), .CLK(clk), .SN(1'b1), .Q(data_out[2])
         );
  DFFSNQ_X1 data_out_reg_1_ ( .D(n707), .CLK(clk), .SN(1'b1), .Q(data_out[1])
         );
  DFFSNQ_X1 data_out_reg_0_ ( .D(n708), .CLK(clk), .SN(1'b1), .Q(data_out[0])
         );
  AND2_X1 U1528 ( .A1(n1736), .A2(n1043), .Z(n979) );
  AND2_X1 U1529 ( .A1(n1198), .A2(n1199), .Z(n1129) );
  OR4_X1 U1530 ( .A1(wr_ptr[40]), .A2(wr_ptr[41]), .A3(wr_ptr[3]), .A4(n1204), 
        .Z(n1201) );
  OR4_X1 U1531 ( .A1(wr_ptr[45]), .A2(wr_ptr[44]), .A3(wr_ptr[43]), .A4(
        wr_ptr[42]), .Z(n1204) );
  OR4_X1 U1532 ( .A1(wr_ptr[17]), .A2(wr_ptr[18]), .A3(wr_ptr[19]), .A4(
        wr_ptr[20]), .Z(n1212) );
  OR4_X1 U1533 ( .A1(wr_ptr[21]), .A2(wr_ptr[22]), .A3(wr_ptr[23]), .A4(
        wr_ptr[24]), .Z(n1211) );
  AND2_X1 U1534 ( .A1(n1335), .A2(n1736), .Z(n1362) );
  XOR2_X1 U1535 ( .A1(n874), .A2(nxt_wr_ptr[51]), .Z(n1374) );
  XOR2_X1 U1536 ( .A1(n872), .A2(nxt_wr_ptr[50]), .Z(n1373) );
  XOR2_X1 U1537 ( .A1(n870), .A2(nxt_wr_ptr[49]), .Z(n1372) );
  XOR2_X1 U1538 ( .A1(n868), .A2(nxt_wr_ptr[48]), .Z(n1371) );
  XOR2_X1 U1539 ( .A1(n882), .A2(nxt_wr_ptr[55]), .Z(n1378) );
  XOR2_X1 U1540 ( .A1(n880), .A2(nxt_wr_ptr[54]), .Z(n1377) );
  XOR2_X1 U1541 ( .A1(n878), .A2(nxt_wr_ptr[53]), .Z(n1376) );
  XOR2_X1 U1542 ( .A1(n876), .A2(nxt_wr_ptr[52]), .Z(n1375) );
  XOR2_X1 U1543 ( .A1(n890), .A2(nxt_wr_ptr[59]), .Z(n1382) );
  XOR2_X1 U1544 ( .A1(n888), .A2(nxt_wr_ptr[58]), .Z(n1381) );
  XOR2_X1 U1545 ( .A1(n886), .A2(nxt_wr_ptr[57]), .Z(n1380) );
  XOR2_X1 U1546 ( .A1(n884), .A2(nxt_wr_ptr[56]), .Z(n1379) );
  XOR2_X1 U1547 ( .A1(n775), .A2(nxt_wr_ptr[63]), .Z(n1386) );
  XOR2_X1 U1548 ( .A1(n896), .A2(nxt_wr_ptr[62]), .Z(n1385) );
  XOR2_X1 U1549 ( .A1(n894), .A2(nxt_wr_ptr[61]), .Z(n1384) );
  XOR2_X1 U1550 ( .A1(n892), .A2(nxt_wr_ptr[60]), .Z(n1383) );
  XOR2_X1 U1551 ( .A1(n842), .A2(nxt_wr_ptr[35]), .Z(n1394) );
  XOR2_X1 U1552 ( .A1(n840), .A2(nxt_wr_ptr[34]), .Z(n1393) );
  XOR2_X1 U1553 ( .A1(n838), .A2(nxt_wr_ptr[33]), .Z(n1392) );
  XOR2_X1 U1554 ( .A1(n836), .A2(nxt_wr_ptr[32]), .Z(n1391) );
  XOR2_X1 U1555 ( .A1(n850), .A2(nxt_wr_ptr[39]), .Z(n1398) );
  XOR2_X1 U1556 ( .A1(n848), .A2(nxt_wr_ptr[38]), .Z(n1397) );
  XOR2_X1 U1557 ( .A1(n846), .A2(nxt_wr_ptr[37]), .Z(n1396) );
  XOR2_X1 U1558 ( .A1(n844), .A2(nxt_wr_ptr[36]), .Z(n1395) );
  XOR2_X1 U1559 ( .A1(n858), .A2(nxt_wr_ptr[43]), .Z(n1402) );
  XOR2_X1 U1560 ( .A1(n856), .A2(nxt_wr_ptr[42]), .Z(n1401) );
  XOR2_X1 U1561 ( .A1(n854), .A2(nxt_wr_ptr[41]), .Z(n1400) );
  XOR2_X1 U1562 ( .A1(n852), .A2(nxt_wr_ptr[40]), .Z(n1399) );
  XOR2_X1 U1563 ( .A1(n866), .A2(nxt_wr_ptr[47]), .Z(n1406) );
  XOR2_X1 U1564 ( .A1(n864), .A2(nxt_wr_ptr[46]), .Z(n1405) );
  XOR2_X1 U1565 ( .A1(n862), .A2(nxt_wr_ptr[45]), .Z(n1404) );
  XOR2_X1 U1566 ( .A1(n860), .A2(nxt_wr_ptr[44]), .Z(n1403) );
  XOR2_X1 U1567 ( .A1(n810), .A2(nxt_wr_ptr[19]), .Z(n1414) );
  XOR2_X1 U1568 ( .A1(n808), .A2(nxt_wr_ptr[18]), .Z(n1413) );
  XOR2_X1 U1569 ( .A1(n806), .A2(nxt_wr_ptr[17]), .Z(n1412) );
  XOR2_X1 U1570 ( .A1(n804), .A2(nxt_wr_ptr[16]), .Z(n1411) );
  XOR2_X1 U1571 ( .A1(n818), .A2(nxt_wr_ptr[23]), .Z(n1418) );
  XOR2_X1 U1572 ( .A1(n816), .A2(nxt_wr_ptr[22]), .Z(n1417) );
  XOR2_X1 U1573 ( .A1(n814), .A2(nxt_wr_ptr[21]), .Z(n1416) );
  XOR2_X1 U1574 ( .A1(n812), .A2(nxt_wr_ptr[20]), .Z(n1415) );
  XOR2_X1 U1575 ( .A1(n826), .A2(nxt_wr_ptr[27]), .Z(n1422) );
  XOR2_X1 U1576 ( .A1(n824), .A2(nxt_wr_ptr[26]), .Z(n1421) );
  XOR2_X1 U1577 ( .A1(n822), .A2(nxt_wr_ptr[25]), .Z(n1420) );
  XOR2_X1 U1578 ( .A1(n820), .A2(nxt_wr_ptr[24]), .Z(n1419) );
  XOR2_X1 U1579 ( .A1(n834), .A2(nxt_wr_ptr[31]), .Z(n1426) );
  XOR2_X1 U1580 ( .A1(n832), .A2(nxt_wr_ptr[30]), .Z(n1425) );
  XOR2_X1 U1581 ( .A1(n830), .A2(nxt_wr_ptr[29]), .Z(n1424) );
  XOR2_X1 U1582 ( .A1(n828), .A2(nxt_wr_ptr[28]), .Z(n1423) );
  XOR2_X1 U1583 ( .A1(n778), .A2(nxt_wr_ptr[3]), .Z(n1434) );
  XOR2_X1 U1584 ( .A1(n777), .A2(nxt_wr_ptr[2]), .Z(n1433) );
  XOR2_X1 U1585 ( .A1(n776), .A2(nxt_wr_ptr[1]), .Z(n1432) );
  XOR2_X1 U1586 ( .A1(n774), .A2(nxt_wr_ptr[0]), .Z(n1431) );
  XOR2_X1 U1587 ( .A1(n786), .A2(nxt_wr_ptr[7]), .Z(n1438) );
  XOR2_X1 U1588 ( .A1(n784), .A2(nxt_wr_ptr[6]), .Z(n1437) );
  XOR2_X1 U1589 ( .A1(n782), .A2(nxt_wr_ptr[5]), .Z(n1436) );
  XOR2_X1 U1590 ( .A1(n780), .A2(nxt_wr_ptr[4]), .Z(n1435) );
  XOR2_X1 U1591 ( .A1(n794), .A2(nxt_wr_ptr[11]), .Z(n1442) );
  XOR2_X1 U1592 ( .A1(n792), .A2(nxt_wr_ptr[10]), .Z(n1441) );
  XOR2_X1 U1593 ( .A1(n790), .A2(nxt_wr_ptr[9]), .Z(n1440) );
  XOR2_X1 U1594 ( .A1(n788), .A2(nxt_wr_ptr[8]), .Z(n1439) );
  XOR2_X1 U1595 ( .A1(n802), .A2(nxt_wr_ptr[15]), .Z(n1446) );
  XOR2_X1 U1596 ( .A1(n800), .A2(nxt_wr_ptr[14]), .Z(n1445) );
  XOR2_X1 U1597 ( .A1(n798), .A2(nxt_wr_ptr[13]), .Z(n1444) );
  XOR2_X1 U1598 ( .A1(n796), .A2(nxt_wr_ptr[12]), .Z(n1443) );
  AND2_X1 U1599 ( .A1(n471), .A2(n1448), .Z(n1273) );
  OR4_X1 U1600 ( .A1(nxt_wr_ptr[53]), .A2(nxt_wr_ptr[54]), .A3(nxt_wr_ptr[55]), 
        .A4(nxt_wr_ptr[56]), .Z(n1457) );
  OR4_X1 U1601 ( .A1(nxt_wr_ptr[57]), .A2(nxt_wr_ptr[58]), .A3(nxt_wr_ptr[59]), 
        .A4(nxt_wr_ptr[5]), .Z(n1456) );
  OR4_X1 U1602 ( .A1(nxt_wr_ptr[60]), .A2(nxt_wr_ptr[61]), .A3(nxt_wr_ptr[62]), 
        .A4(nxt_wr_ptr[63]), .Z(n1455) );
  OR4_X1 U1603 ( .A1(nxt_wr_ptr[6]), .A2(nxt_wr_ptr[7]), .A3(nxt_wr_ptr[8]), 
        .A4(nxt_wr_ptr[9]), .Z(n1454) );
  OR4_X1 U1604 ( .A1(nxt_wr_ptr[39]), .A2(nxt_wr_ptr[3]), .A3(nxt_wr_ptr[40]), 
        .A4(nxt_wr_ptr[41]), .Z(n1461) );
  OR4_X1 U1605 ( .A1(nxt_wr_ptr[42]), .A2(nxt_wr_ptr[43]), .A3(nxt_wr_ptr[44]), 
        .A4(nxt_wr_ptr[45]), .Z(n1460) );
  OR4_X1 U1606 ( .A1(nxt_wr_ptr[24]), .A2(nxt_wr_ptr[25]), .A3(nxt_wr_ptr[26]), 
        .A4(nxt_wr_ptr[27]), .Z(n1465) );
  OR4_X1 U1607 ( .A1(nxt_wr_ptr[28]), .A2(nxt_wr_ptr[29]), .A3(nxt_wr_ptr[2]), 
        .A4(nxt_wr_ptr[30]), .Z(n1464) );
  OR4_X1 U1608 ( .A1(nxt_wr_ptr[31]), .A2(nxt_wr_ptr[32]), .A3(nxt_wr_ptr[33]), 
        .A4(nxt_wr_ptr[34]), .Z(n1463) );
  OR4_X1 U1609 ( .A1(nxt_wr_ptr[35]), .A2(nxt_wr_ptr[36]), .A3(nxt_wr_ptr[37]), 
        .A4(nxt_wr_ptr[38]), .Z(n1462) );
  OR4_X1 U1610 ( .A1(nxt_wr_ptr[13]), .A2(nxt_wr_ptr[14]), .A3(nxt_wr_ptr[15]), 
        .A4(nxt_wr_ptr[16]), .Z(n1468) );
  OR4_X1 U1611 ( .A1(nxt_wr_ptr[17]), .A2(nxt_wr_ptr[18]), .A3(nxt_wr_ptr[19]), 
        .A4(nxt_wr_ptr[1]), .Z(n1467) );
  OR4_X1 U1612 ( .A1(nxt_wr_ptr[20]), .A2(nxt_wr_ptr[21]), .A3(nxt_wr_ptr[22]), 
        .A4(nxt_wr_ptr[23]), .Z(n1466) );
  AND2_X1 U1613 ( .A1(wr), .A2(n1712), .Z(n1130) );
  circ_q_WORD_SZ64_1_DW01_inc_0 add_97 ( .A(nxt_wr_ptr), .SUM({N595, N594, 
        N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, 
        N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, 
        N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, 
        N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, 
        N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, 
        N533, N532}) );
  circ_q_WORD_SZ64_1_DW01_inc_1 add_72 ( .A(nxt_rd_ptr), .SUM({N309, N308, 
        N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, 
        N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, 
        N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, 
        N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, 
        N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, 
        N247, N246}) );
  BUF_X2 U4 ( .I(n950), .Z(n471) );
  BUF_X2 U452 ( .I(n1273), .Z(n484) );
  BUF_X2 U453 ( .I(n1273), .Z(n483) );
  BUF_X2 U454 ( .I(n1273), .Z(n479) );
  BUF_X2 U455 ( .I(n1273), .Z(n480) );
  BUF_X2 U456 ( .I(n1273), .Z(n481) );
  BUF_X2 U457 ( .I(n1273), .Z(n482) );
  BUF_X2 U458 ( .I(n1339), .Z(n477) );
  BUF_X2 U459 ( .I(n1339), .Z(n472) );
  BUF_X2 U460 ( .I(n1339), .Z(n473) );
  BUF_X2 U461 ( .I(n1339), .Z(n474) );
  BUF_X2 U462 ( .I(n1339), .Z(n475) );
  BUF_X2 U463 ( .I(n1339), .Z(n476) );
  BUF_X2 U464 ( .I(n950), .Z(n470) );
  BUF_X2 U465 ( .I(n950), .Z(n469) );
  BUF_X2 U466 ( .I(n950), .Z(n468) );
  BUF_X2 U467 ( .I(n950), .Z(n467) );
  INV_X1 U468 ( .I(n564), .ZN(n532) );
  INV_X1 U469 ( .I(n564), .ZN(n533) );
  INV_X1 U470 ( .I(n564), .ZN(n534) );
  INV_X1 U471 ( .I(n515), .ZN(n524) );
  INV_X1 U472 ( .I(n565), .ZN(n535) );
  INV_X1 U473 ( .I(n565), .ZN(n536) );
  INV_X1 U474 ( .I(n456), .ZN(n950) );
  NAND2_X1 U475 ( .A1(n449), .A2(n1341), .ZN(n1339) );
  BUF_X2 U476 ( .I(n709), .Z(n462) );
  BUF_X2 U477 ( .I(n979), .Z(n571) );
  BUF_X2 U478 ( .I(n578), .Z(n577) );
  BUF_X2 U479 ( .I(n579), .Z(n573) );
  BUF_X2 U480 ( .I(n579), .Z(n574) );
  BUF_X2 U481 ( .I(n579), .Z(n572) );
  BUF_X2 U482 ( .I(n578), .Z(n575) );
  BUF_X2 U483 ( .I(n578), .Z(n576) );
  INV_X1 U484 ( .I(n449), .ZN(n478) );
  BUF_X2 U485 ( .I(n516), .Z(n515) );
  BUF_X2 U486 ( .I(n979), .Z(n570) );
  BUF_X2 U487 ( .I(n979), .Z(n566) );
  BUF_X2 U488 ( .I(n979), .Z(n567) );
  BUF_X2 U489 ( .I(n979), .Z(n568) );
  BUF_X2 U490 ( .I(n979), .Z(n569) );
  INV_X1 U491 ( .I(n493), .ZN(n487) );
  INV_X1 U492 ( .I(n493), .ZN(n489) );
  INV_X1 U493 ( .I(n493), .ZN(n488) );
  BUF_X2 U494 ( .I(n709), .Z(n465) );
  BUF_X2 U495 ( .I(n709), .Z(n464) );
  BUF_X2 U496 ( .I(n709), .Z(n463) );
  BUF_X2 U497 ( .I(n709), .Z(n461) );
  BUF_X2 U498 ( .I(n709), .Z(n460) );
  BUF_X2 U499 ( .I(n709), .Z(n459) );
  BUF_X2 U500 ( .I(n709), .Z(n458) );
  BUF_X2 U501 ( .I(n709), .Z(n457) );
  BUF_X2 U502 ( .I(n516), .Z(n514) );
  BUF_X2 U503 ( .I(n517), .Z(n513) );
  BUF_X2 U504 ( .I(n517), .Z(n512) );
  BUF_X2 U505 ( .I(n517), .Z(n511) );
  BUF_X2 U506 ( .I(n518), .Z(n510) );
  BUF_X2 U507 ( .I(n518), .Z(n509) );
  BUF_X2 U508 ( .I(n518), .Z(n508) );
  BUF_X2 U509 ( .I(n519), .Z(n507) );
  BUF_X2 U510 ( .I(n519), .Z(n506) );
  BUF_X2 U511 ( .I(n519), .Z(n505) );
  BUF_X2 U512 ( .I(n520), .Z(n504) );
  BUF_X2 U513 ( .I(n520), .Z(n503) );
  BUF_X2 U514 ( .I(n520), .Z(n502) );
  BUF_X2 U515 ( .I(n521), .Z(n501) );
  BUF_X2 U516 ( .I(n521), .Z(n500) );
  BUF_X2 U517 ( .I(n521), .Z(n499) );
  BUF_X2 U518 ( .I(n522), .Z(n498) );
  BUF_X2 U519 ( .I(n522), .Z(n497) );
  BUF_X2 U520 ( .I(n522), .Z(n496) );
  BUF_X2 U521 ( .I(n523), .Z(n495) );
  BUF_X2 U522 ( .I(n523), .Z(n494) );
  BUF_X2 U523 ( .I(n709), .Z(n466) );
  INV_X1 U524 ( .I(n492), .ZN(n485) );
  INV_X1 U525 ( .I(n491), .ZN(n486) );
  OAI22_X1 U526 ( .A1(n896), .A2(n462), .B1(n472), .B2(n712), .ZN(n1545) );
  INV_X1 U527 ( .I(N308), .ZN(n712) );
  OAI22_X1 U528 ( .A1(n894), .A2(n462), .B1(n472), .B2(n713), .ZN(n1546) );
  INV_X1 U529 ( .I(N307), .ZN(n713) );
  OAI22_X1 U530 ( .A1(n892), .A2(n462), .B1(n472), .B2(n714), .ZN(n1547) );
  INV_X1 U531 ( .I(N306), .ZN(n714) );
  OAI22_X1 U532 ( .A1(n890), .A2(n462), .B1(n472), .B2(n715), .ZN(n1548) );
  INV_X1 U533 ( .I(N305), .ZN(n715) );
  OAI22_X1 U534 ( .A1(n888), .A2(n461), .B1(n472), .B2(n716), .ZN(n1549) );
  INV_X1 U535 ( .I(N304), .ZN(n716) );
  OAI22_X1 U536 ( .A1(n886), .A2(n461), .B1(n472), .B2(n717), .ZN(n1550) );
  INV_X1 U537 ( .I(N303), .ZN(n717) );
  OAI22_X1 U538 ( .A1(n884), .A2(n461), .B1(n472), .B2(n718), .ZN(n1551) );
  INV_X1 U539 ( .I(N302), .ZN(n718) );
  OAI22_X1 U540 ( .A1(n882), .A2(n461), .B1(n472), .B2(n719), .ZN(n1552) );
  INV_X1 U541 ( .I(N301), .ZN(n719) );
  OAI22_X1 U542 ( .A1(n880), .A2(n461), .B1(n472), .B2(n720), .ZN(n1553) );
  INV_X1 U543 ( .I(N300), .ZN(n720) );
  OAI22_X1 U544 ( .A1(n878), .A2(n461), .B1(n472), .B2(n721), .ZN(n1554) );
  INV_X1 U545 ( .I(N299), .ZN(n721) );
  OAI22_X1 U546 ( .A1(n876), .A2(n461), .B1(n472), .B2(n722), .ZN(n1555) );
  INV_X1 U547 ( .I(N298), .ZN(n722) );
  OAI22_X1 U548 ( .A1(n874), .A2(n461), .B1(n472), .B2(n723), .ZN(n1556) );
  INV_X1 U549 ( .I(N297), .ZN(n723) );
  OAI22_X1 U550 ( .A1(n872), .A2(n461), .B1(n473), .B2(n724), .ZN(n1557) );
  INV_X1 U551 ( .I(N296), .ZN(n724) );
  OAI22_X1 U552 ( .A1(n870), .A2(n461), .B1(n473), .B2(n725), .ZN(n1558) );
  INV_X1 U553 ( .I(N295), .ZN(n725) );
  OAI22_X1 U554 ( .A1(n868), .A2(n461), .B1(n473), .B2(n726), .ZN(n1559) );
  INV_X1 U555 ( .I(N294), .ZN(n726) );
  OAI22_X1 U556 ( .A1(n866), .A2(n461), .B1(n473), .B2(n727), .ZN(n1560) );
  INV_X1 U557 ( .I(N293), .ZN(n727) );
  OAI22_X1 U558 ( .A1(n864), .A2(n460), .B1(n473), .B2(n728), .ZN(n1561) );
  INV_X1 U559 ( .I(N292), .ZN(n728) );
  OAI22_X1 U560 ( .A1(n862), .A2(n460), .B1(n473), .B2(n729), .ZN(n1562) );
  INV_X1 U561 ( .I(N291), .ZN(n729) );
  OAI22_X1 U562 ( .A1(n860), .A2(n460), .B1(n473), .B2(n730), .ZN(n1563) );
  INV_X1 U563 ( .I(N290), .ZN(n730) );
  OAI22_X1 U564 ( .A1(n858), .A2(n460), .B1(n473), .B2(n731), .ZN(n1564) );
  INV_X1 U565 ( .I(N289), .ZN(n731) );
  OAI22_X1 U566 ( .A1(n856), .A2(n460), .B1(n473), .B2(n732), .ZN(n1565) );
  INV_X1 U567 ( .I(N288), .ZN(n732) );
  OAI22_X1 U568 ( .A1(n854), .A2(n460), .B1(n473), .B2(n733), .ZN(n1566) );
  INV_X1 U569 ( .I(N287), .ZN(n733) );
  OAI22_X1 U570 ( .A1(n852), .A2(n460), .B1(n473), .B2(n734), .ZN(n1567) );
  INV_X1 U571 ( .I(N286), .ZN(n734) );
  OAI22_X1 U572 ( .A1(n850), .A2(n460), .B1(n473), .B2(n735), .ZN(n1568) );
  INV_X1 U573 ( .I(N285), .ZN(n735) );
  OAI22_X1 U574 ( .A1(n848), .A2(n460), .B1(n474), .B2(n736), .ZN(n1569) );
  INV_X1 U575 ( .I(N284), .ZN(n736) );
  OAI22_X1 U576 ( .A1(n846), .A2(n460), .B1(n474), .B2(n737), .ZN(n1570) );
  INV_X1 U577 ( .I(N283), .ZN(n737) );
  OAI22_X1 U578 ( .A1(n844), .A2(n460), .B1(n474), .B2(n738), .ZN(n1571) );
  INV_X1 U579 ( .I(N282), .ZN(n738) );
  OAI22_X1 U580 ( .A1(n842), .A2(n460), .B1(n474), .B2(n739), .ZN(n1572) );
  INV_X1 U581 ( .I(N281), .ZN(n739) );
  OAI22_X1 U582 ( .A1(n840), .A2(n459), .B1(n474), .B2(n740), .ZN(n1573) );
  INV_X1 U583 ( .I(N280), .ZN(n740) );
  OAI22_X1 U584 ( .A1(n838), .A2(n459), .B1(n474), .B2(n741), .ZN(n1574) );
  INV_X1 U585 ( .I(N279), .ZN(n741) );
  OAI22_X1 U586 ( .A1(n836), .A2(n459), .B1(n474), .B2(n742), .ZN(n1575) );
  INV_X1 U587 ( .I(N278), .ZN(n742) );
  OAI22_X1 U588 ( .A1(n834), .A2(n459), .B1(n474), .B2(n743), .ZN(n1576) );
  INV_X1 U589 ( .I(N277), .ZN(n743) );
  OAI22_X1 U590 ( .A1(n832), .A2(n459), .B1(n474), .B2(n744), .ZN(n1577) );
  INV_X1 U591 ( .I(N276), .ZN(n744) );
  OAI22_X1 U592 ( .A1(n830), .A2(n459), .B1(n474), .B2(n745), .ZN(n1578) );
  INV_X1 U593 ( .I(N275), .ZN(n745) );
  OAI22_X1 U594 ( .A1(n828), .A2(n459), .B1(n474), .B2(n746), .ZN(n1579) );
  INV_X1 U595 ( .I(N274), .ZN(n746) );
  OAI22_X1 U596 ( .A1(n826), .A2(n459), .B1(n474), .B2(n747), .ZN(n1580) );
  INV_X1 U597 ( .I(N273), .ZN(n747) );
  OAI22_X1 U598 ( .A1(n824), .A2(n459), .B1(n475), .B2(n748), .ZN(n1581) );
  INV_X1 U599 ( .I(N272), .ZN(n748) );
  OAI22_X1 U600 ( .A1(n822), .A2(n459), .B1(n475), .B2(n749), .ZN(n1582) );
  INV_X1 U601 ( .I(N271), .ZN(n749) );
  OAI22_X1 U602 ( .A1(n820), .A2(n459), .B1(n475), .B2(n750), .ZN(n1583) );
  INV_X1 U603 ( .I(N270), .ZN(n750) );
  OAI22_X1 U604 ( .A1(n818), .A2(n459), .B1(n475), .B2(n751), .ZN(n1584) );
  INV_X1 U605 ( .I(N269), .ZN(n751) );
  OAI22_X1 U606 ( .A1(n816), .A2(n458), .B1(n475), .B2(n752), .ZN(n1585) );
  INV_X1 U607 ( .I(N268), .ZN(n752) );
  OAI22_X1 U608 ( .A1(n814), .A2(n458), .B1(n475), .B2(n753), .ZN(n1586) );
  INV_X1 U609 ( .I(N267), .ZN(n753) );
  OAI22_X1 U610 ( .A1(n812), .A2(n458), .B1(n475), .B2(n754), .ZN(n1587) );
  INV_X1 U611 ( .I(N266), .ZN(n754) );
  OAI22_X1 U612 ( .A1(n810), .A2(n458), .B1(n475), .B2(n755), .ZN(n1588) );
  INV_X1 U613 ( .I(N265), .ZN(n755) );
  OAI22_X1 U614 ( .A1(n808), .A2(n458), .B1(n475), .B2(n756), .ZN(n1589) );
  INV_X1 U615 ( .I(N264), .ZN(n756) );
  OAI22_X1 U616 ( .A1(n806), .A2(n458), .B1(n475), .B2(n757), .ZN(n1590) );
  INV_X1 U617 ( .I(N263), .ZN(n757) );
  OAI22_X1 U618 ( .A1(n804), .A2(n458), .B1(n475), .B2(n758), .ZN(n1591) );
  INV_X1 U619 ( .I(N262), .ZN(n758) );
  INV_X1 U620 ( .I(n1219), .ZN(n490) );
  BUF_X2 U621 ( .I(n1230), .Z(n456) );
  NAND2_X1 U622 ( .A1(n490), .A2(n1736), .ZN(n1230) );
  OAI22_X1 U623 ( .A1(n802), .A2(n458), .B1(n475), .B2(n759), .ZN(n1592) );
  INV_X1 U624 ( .I(N261), .ZN(n759) );
  INV_X1 U625 ( .I(n1338), .ZN(n709) );
  AND2_X1 U626 ( .A1(n462), .A2(n1736), .Z(n449) );
  OAI22_X1 U627 ( .A1(n777), .A2(n457), .B1(n477), .B2(n772), .ZN(n1605) );
  INV_X1 U628 ( .I(N248), .ZN(n772) );
  OAI22_X1 U629 ( .A1(n776), .A2(n457), .B1(n477), .B2(n773), .ZN(n1606) );
  INV_X1 U630 ( .I(N247), .ZN(n773) );
  OAI22_X1 U631 ( .A1(n800), .A2(n458), .B1(n476), .B2(n760), .ZN(n1593) );
  INV_X1 U632 ( .I(N260), .ZN(n760) );
  OAI22_X1 U633 ( .A1(n798), .A2(n458), .B1(n476), .B2(n761), .ZN(n1594) );
  INV_X1 U634 ( .I(N259), .ZN(n761) );
  OAI22_X1 U635 ( .A1(n796), .A2(n458), .B1(n476), .B2(n762), .ZN(n1595) );
  INV_X1 U636 ( .I(N258), .ZN(n762) );
  OAI22_X1 U637 ( .A1(n794), .A2(n458), .B1(n476), .B2(n763), .ZN(n1596) );
  INV_X1 U638 ( .I(N257), .ZN(n763) );
  OAI22_X1 U639 ( .A1(n792), .A2(n457), .B1(n476), .B2(n764), .ZN(n1597) );
  INV_X1 U640 ( .I(N256), .ZN(n764) );
  OAI22_X1 U641 ( .A1(n790), .A2(n457), .B1(n476), .B2(n765), .ZN(n1598) );
  INV_X1 U642 ( .I(N255), .ZN(n765) );
  OAI22_X1 U643 ( .A1(n788), .A2(n457), .B1(n476), .B2(n766), .ZN(n1599) );
  INV_X1 U644 ( .I(N254), .ZN(n766) );
  OAI22_X1 U645 ( .A1(n786), .A2(n457), .B1(n476), .B2(n767), .ZN(n1600) );
  INV_X1 U646 ( .I(N253), .ZN(n767) );
  OAI22_X1 U647 ( .A1(n784), .A2(n457), .B1(n476), .B2(n768), .ZN(n1601) );
  INV_X1 U648 ( .I(N252), .ZN(n768) );
  OAI22_X1 U649 ( .A1(n782), .A2(n457), .B1(n476), .B2(n769), .ZN(n1602) );
  INV_X1 U650 ( .I(N251), .ZN(n769) );
  OAI22_X1 U651 ( .A1(n780), .A2(n457), .B1(n476), .B2(n770), .ZN(n1603) );
  INV_X1 U652 ( .I(N250), .ZN(n770) );
  OAI22_X1 U653 ( .A1(n778), .A2(n457), .B1(n476), .B2(n771), .ZN(n1604) );
  INV_X1 U654 ( .I(N249), .ZN(n771) );
  NAND4_X1 U655 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043)
         );
  NOR4_X1 U656 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1044) );
  NOR4_X1 U657 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1045) );
  BUF_X2 U658 ( .I(n978), .Z(n579) );
  BUF_X2 U659 ( .I(n978), .Z(n578) );
  OAI22_X1 U660 ( .A1(n462), .A2(n779), .B1(n778), .B2(n478), .ZN(n1543) );
  OAI22_X1 U661 ( .A1(n464), .A2(n851), .B1(n850), .B2(n478), .ZN(n1507) );
  OAI22_X1 U662 ( .A1(n464), .A2(n849), .B1(n848), .B2(n478), .ZN(n1508) );
  OAI22_X1 U663 ( .A1(n464), .A2(n847), .B1(n846), .B2(n478), .ZN(n1509) );
  OAI22_X1 U664 ( .A1(n464), .A2(n845), .B1(n844), .B2(n478), .ZN(n1510) );
  OAI22_X1 U665 ( .A1(n464), .A2(n843), .B1(n842), .B2(n478), .ZN(n1511) );
  OAI22_X1 U666 ( .A1(n464), .A2(n841), .B1(n840), .B2(n478), .ZN(n1512) );
  OAI22_X1 U667 ( .A1(n464), .A2(n839), .B1(n838), .B2(n478), .ZN(n1513) );
  OAI22_X1 U668 ( .A1(n464), .A2(n837), .B1(n836), .B2(n478), .ZN(n1514) );
  OAI22_X1 U669 ( .A1(n464), .A2(n835), .B1(n834), .B2(n478), .ZN(n1515) );
  OAI22_X1 U670 ( .A1(n464), .A2(n833), .B1(n832), .B2(n478), .ZN(n1516) );
  OAI22_X1 U671 ( .A1(n464), .A2(n831), .B1(n830), .B2(n478), .ZN(n1517) );
  OAI22_X1 U672 ( .A1(n464), .A2(n829), .B1(n828), .B2(n478), .ZN(n1518) );
  OAI22_X1 U673 ( .A1(n464), .A2(n827), .B1(n826), .B2(n478), .ZN(n1519) );
  OAI22_X1 U674 ( .A1(n464), .A2(n825), .B1(n824), .B2(n478), .ZN(n1520) );
  OAI22_X1 U675 ( .A1(n463), .A2(n823), .B1(n822), .B2(n478), .ZN(n1521) );
  OAI22_X1 U676 ( .A1(n463), .A2(n821), .B1(n820), .B2(n478), .ZN(n1522) );
  OAI22_X1 U677 ( .A1(n463), .A2(n819), .B1(n818), .B2(n478), .ZN(n1523) );
  OAI22_X1 U678 ( .A1(n463), .A2(n817), .B1(n816), .B2(n478), .ZN(n1524) );
  OAI22_X1 U679 ( .A1(n463), .A2(n815), .B1(n814), .B2(n478), .ZN(n1525) );
  OAI22_X1 U680 ( .A1(n463), .A2(n813), .B1(n812), .B2(n478), .ZN(n1526) );
  OAI22_X1 U681 ( .A1(n463), .A2(n811), .B1(n810), .B2(n478), .ZN(n1527) );
  OAI22_X1 U682 ( .A1(n463), .A2(n809), .B1(n808), .B2(n478), .ZN(n1528) );
  OAI22_X1 U683 ( .A1(n463), .A2(n807), .B1(n806), .B2(n478), .ZN(n1529) );
  OAI22_X1 U684 ( .A1(n463), .A2(n805), .B1(n804), .B2(n478), .ZN(n1530) );
  OAI22_X1 U685 ( .A1(n463), .A2(n803), .B1(n802), .B2(n478), .ZN(n1531) );
  OAI22_X1 U686 ( .A1(n463), .A2(n801), .B1(n800), .B2(n478), .ZN(n1532) );
  OAI22_X1 U687 ( .A1(n463), .A2(n799), .B1(n798), .B2(n478), .ZN(n1533) );
  OAI22_X1 U688 ( .A1(n463), .A2(n797), .B1(n796), .B2(n478), .ZN(n1534) );
  OAI22_X1 U689 ( .A1(n462), .A2(n795), .B1(n794), .B2(n478), .ZN(n1535) );
  OAI22_X1 U690 ( .A1(n462), .A2(n793), .B1(n792), .B2(n478), .ZN(n1536) );
  OAI22_X1 U691 ( .A1(n462), .A2(n791), .B1(n790), .B2(n478), .ZN(n1537) );
  OAI22_X1 U692 ( .A1(n462), .A2(n789), .B1(n788), .B2(n478), .ZN(n1538) );
  OAI22_X1 U693 ( .A1(n462), .A2(n787), .B1(n786), .B2(n478), .ZN(n1539) );
  OAI22_X1 U694 ( .A1(n462), .A2(n785), .B1(n784), .B2(n478), .ZN(n1540) );
  OAI22_X1 U695 ( .A1(n462), .A2(n783), .B1(n782), .B2(n478), .ZN(n1541) );
  OAI22_X1 U696 ( .A1(n462), .A2(n781), .B1(n780), .B2(n478), .ZN(n1542) );
  OAI22_X1 U697 ( .A1(n466), .A2(n893), .B1(n892), .B2(n478), .ZN(n1486) );
  OAI22_X1 U698 ( .A1(n466), .A2(n887), .B1(n886), .B2(n478), .ZN(n1489) );
  OAI22_X1 U699 ( .A1(n465), .A2(n879), .B1(n878), .B2(n478), .ZN(n1493) );
  OAI22_X1 U700 ( .A1(n465), .A2(n865), .B1(n864), .B2(n478), .ZN(n1500) );
  OAI22_X1 U701 ( .A1(n465), .A2(n857), .B1(n856), .B2(n478), .ZN(n1504) );
  OAI22_X1 U702 ( .A1(n466), .A2(n898), .B1(n775), .B2(n478), .ZN(n1483) );
  OAI22_X1 U703 ( .A1(n466), .A2(n895), .B1(n894), .B2(n478), .ZN(n1485) );
  OAI22_X1 U704 ( .A1(n466), .A2(n889), .B1(n888), .B2(n478), .ZN(n1488) );
  OAI22_X1 U705 ( .A1(n466), .A2(n881), .B1(n880), .B2(n478), .ZN(n1492) );
  OAI22_X1 U706 ( .A1(n465), .A2(n873), .B1(n872), .B2(n478), .ZN(n1496) );
  OAI22_X1 U707 ( .A1(n465), .A2(n867), .B1(n866), .B2(n478), .ZN(n1499) );
  OAI22_X1 U708 ( .A1(n465), .A2(n859), .B1(n858), .B2(n478), .ZN(n1503) );
  OAI22_X1 U709 ( .A1(n466), .A2(n897), .B1(n896), .B2(n478), .ZN(n1484) );
  OAI22_X1 U710 ( .A1(n466), .A2(n891), .B1(n890), .B2(n478), .ZN(n1487) );
  OAI22_X1 U711 ( .A1(n466), .A2(n883), .B1(n882), .B2(n478), .ZN(n1491) );
  OAI22_X1 U712 ( .A1(n465), .A2(n875), .B1(n874), .B2(n478), .ZN(n1495) );
  OAI22_X1 U713 ( .A1(n465), .A2(n869), .B1(n868), .B2(n478), .ZN(n1498) );
  OAI22_X1 U714 ( .A1(n465), .A2(n861), .B1(n860), .B2(n478), .ZN(n1502) );
  OAI22_X1 U715 ( .A1(n465), .A2(n853), .B1(n852), .B2(n478), .ZN(n1506) );
  OAI22_X1 U716 ( .A1(n466), .A2(n885), .B1(n884), .B2(n478), .ZN(n1490) );
  OAI22_X1 U717 ( .A1(n465), .A2(n877), .B1(n876), .B2(n478), .ZN(n1494) );
  OAI22_X1 U718 ( .A1(n465), .A2(n871), .B1(n870), .B2(n478), .ZN(n1497) );
  OAI22_X1 U719 ( .A1(n465), .A2(n863), .B1(n862), .B2(n478), .ZN(n1501) );
  OAI22_X1 U720 ( .A1(n465), .A2(n855), .B1(n854), .B2(n478), .ZN(n1505) );
  BUF_X2 U721 ( .I(n1065), .Z(n531) );
  BUF_X2 U722 ( .I(n1133), .Z(n516) );
  INV_X1 U723 ( .I(n1219), .ZN(n493) );
  NOR4_X1 U724 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
  NAND4_X1 U725 ( .A1(n785), .A2(n787), .A3(n789), .A4(n791), .ZN(n1048) );
  NAND4_X1 U726 ( .A1(n893), .A2(n895), .A3(n897), .A4(n898), .ZN(n1049) );
  NAND4_X1 U727 ( .A1(n887), .A2(n889), .A3(n891), .A4(n783), .ZN(n1050) );
  NAND4_X1 U728 ( .A1(n879), .A2(n881), .A3(n883), .A4(n885), .ZN(n1051) );
  NOR4_X1 U729 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1046) );
  NAND4_X1 U730 ( .A1(n781), .A2(n873), .A3(n875), .A4(n877), .ZN(n1052) );
  NAND4_X1 U731 ( .A1(n865), .A2(n867), .A3(n869), .A4(n871), .ZN(n1053) );
  NAND4_X1 U732 ( .A1(n857), .A2(n859), .A3(n861), .A4(n863), .ZN(n1054) );
  NAND4_X1 U733 ( .A1(n851), .A2(n779), .A3(n853), .A4(n855), .ZN(n1055) );
  NAND4_X1 U734 ( .A1(n819), .A2(n821), .A3(n823), .A4(n825), .ZN(n1059) );
  NAND4_X1 U735 ( .A1(n827), .A2(n829), .A3(n831), .A4(n833), .ZN(n1058) );
  NAND4_X1 U736 ( .A1(n795), .A2(n797), .A3(n799), .A4(n801), .ZN(n1062) );
  NAND4_X1 U737 ( .A1(n835), .A2(n837), .A3(n839), .A4(n841), .ZN(n1057) );
  NAND4_X1 U738 ( .A1(n803), .A2(n805), .A3(n807), .A4(n809), .ZN(n1061) );
  NAND4_X1 U739 ( .A1(n843), .A2(n845), .A3(n847), .A4(n849), .ZN(n1056) );
  OAI22_X1 U740 ( .A1(n492), .A2(n1712), .B1(n456), .B2(n1335), .ZN(n1482) );
  OAI22_X1 U741 ( .A1(n490), .A2(n1733), .B1(n456), .B2(n1732), .ZN(n1471) );
  OAI22_X1 U742 ( .A1(n493), .A2(n1735), .B1(n456), .B2(n1734), .ZN(n1470) );
  OAI22_X1 U743 ( .A1(n492), .A2(n1731), .B1(n456), .B2(n1730), .ZN(n1472) );
  OAI22_X1 U744 ( .A1(n491), .A2(n1729), .B1(n456), .B2(n1728), .ZN(n1473) );
  OAI22_X1 U745 ( .A1(n491), .A2(n1727), .B1(n456), .B2(n1726), .ZN(n1474) );
  OAI22_X1 U746 ( .A1(n491), .A2(n1725), .B1(n456), .B2(n1724), .ZN(n1475) );
  OAI22_X1 U747 ( .A1(n492), .A2(n1723), .B1(n456), .B2(n1722), .ZN(n1476) );
  OAI22_X1 U748 ( .A1(n493), .A2(n1721), .B1(n456), .B2(n1720), .ZN(n1477) );
  OAI22_X1 U749 ( .A1(n492), .A2(n1719), .B1(n456), .B2(n1718), .ZN(n1478) );
  OAI22_X1 U750 ( .A1(n492), .A2(n1717), .B1(n456), .B2(n1716), .ZN(n1479) );
  OAI22_X1 U751 ( .A1(n491), .A2(n1715), .B1(n456), .B2(n1714), .ZN(n1480) );
  BUF_X2 U752 ( .I(n1133), .Z(n517) );
  BUF_X2 U753 ( .I(n1133), .Z(n518) );
  BUF_X2 U754 ( .I(n1133), .Z(n519) );
  BUF_X2 U755 ( .I(n1133), .Z(n520) );
  BUF_X2 U756 ( .I(n1133), .Z(n521) );
  BUF_X2 U757 ( .I(n1133), .Z(n522) );
  BUF_X2 U758 ( .I(n1133), .Z(n523) );
  NAND4_X1 U759 ( .A1(n811), .A2(n813), .A3(n815), .A4(n817), .ZN(n1060) );
  INV_X1 U760 ( .I(n1219), .ZN(n491) );
  INV_X1 U761 ( .I(n1219), .ZN(n492) );
  BUF_X2 U762 ( .I(n1065), .Z(n530) );
  BUF_X2 U763 ( .I(n1065), .Z(n529) );
  BUF_X2 U764 ( .I(n1065), .Z(n528) );
  BUF_X2 U765 ( .I(n1065), .Z(n527) );
  BUF_X2 U766 ( .I(n1065), .Z(n526) );
  BUF_X2 U767 ( .I(n1065), .Z(n525) );
  NAND4_X1 U768 ( .A1(n1723), .A2(n1725), .A3(n1727), .A4(n1729), .ZN(n1203)
         );
  NAND4_X1 U769 ( .A1(n1715), .A2(n1731), .A3(n1733), .A4(n1735), .ZN(n1202)
         );
  NAND4_X1 U770 ( .A1(n1450), .A2(n1451), .A3(n1452), .A4(n1453), .ZN(n1448)
         );
  NOR4_X1 U771 ( .A1(n1466), .A2(n1467), .A3(n1468), .A4(n1469), .ZN(n1450) );
  NOR4_X1 U772 ( .A1(n1462), .A2(n1463), .A3(n1464), .A4(n1465), .ZN(n1451) );
  NOR4_X1 U773 ( .A1(n1458), .A2(n1459), .A3(n1460), .A4(n1461), .ZN(n1452) );
  NAND4_X1 U774 ( .A1(n1722), .A2(n1724), .A3(n1726), .A4(n1728), .ZN(n1459)
         );
  NAND4_X1 U775 ( .A1(n1714), .A2(n1730), .A3(n1732), .A4(n1734), .ZN(n1458)
         );
  OAI21_X1 U776 ( .A1(n1338), .A2(n1362), .B(n710), .ZN(n1609) );
  NAND4_X1 U777 ( .A1(n1342), .A2(n1343), .A3(n1344), .A4(n1345), .ZN(n1341)
         );
  NOR4_X1 U778 ( .A1(n1358), .A2(n1359), .A3(n1360), .A4(n1361), .ZN(n1342) );
  NOR4_X1 U779 ( .A1(n1354), .A2(n1355), .A3(n1356), .A4(n1357), .ZN(n1343) );
  NOR4_X1 U780 ( .A1(n1350), .A2(n1351), .A3(n1352), .A4(n1353), .ZN(n1344) );
  NOR4_X1 U781 ( .A1(n1346), .A2(n1347), .A3(n1348), .A4(n1349), .ZN(n1345) );
  NAND4_X1 U782 ( .A1(n784), .A2(n786), .A3(n788), .A4(n790), .ZN(n1346) );
  NAND4_X1 U783 ( .A1(n886), .A2(n888), .A3(n890), .A4(n782), .ZN(n1348) );
  NAND4_X1 U784 ( .A1(n878), .A2(n880), .A3(n882), .A4(n884), .ZN(n1349) );
  NAND4_X1 U785 ( .A1(n850), .A2(n778), .A3(n852), .A4(n854), .ZN(n1353) );
  NAND4_X1 U786 ( .A1(n892), .A2(n894), .A3(n896), .A4(n775), .ZN(n1347) );
  NAND4_X1 U787 ( .A1(n820), .A2(n822), .A3(n824), .A4(n826), .ZN(n1357) );
  NAND4_X1 U788 ( .A1(n856), .A2(n858), .A3(n860), .A4(n862), .ZN(n1352) );
  NAND4_X1 U789 ( .A1(n828), .A2(n830), .A3(n777), .A4(n832), .ZN(n1356) );
  NAND4_X1 U790 ( .A1(n864), .A2(n866), .A3(n868), .A4(n870), .ZN(n1351) );
  NAND4_X1 U791 ( .A1(n834), .A2(n836), .A3(n838), .A4(n840), .ZN(n1355) );
  NAND4_X1 U792 ( .A1(n798), .A2(n800), .A3(n802), .A4(n804), .ZN(n1360) );
  NAND4_X1 U793 ( .A1(n806), .A2(n808), .A3(n810), .A4(n776), .ZN(n1359) );
  NAND4_X1 U794 ( .A1(n780), .A2(n872), .A3(n874), .A4(n876), .ZN(n1350) );
  NAND4_X1 U795 ( .A1(n842), .A2(n844), .A3(n846), .A4(n848), .ZN(n1354) );
  NAND4_X1 U796 ( .A1(n812), .A2(n814), .A3(n816), .A4(n818), .ZN(n1358) );
  NAND4_X1 U797 ( .A1(n1363), .A2(n1364), .A3(n1365), .A4(n1366), .ZN(n1335)
         );
  NOR4_X1 U798 ( .A1(n1407), .A2(n1408), .A3(n1409), .A4(n1410), .ZN(n1364) );
  NOR4_X1 U799 ( .A1(n1387), .A2(n1388), .A3(n1389), .A4(n1390), .ZN(n1365) );
  NOR4_X1 U800 ( .A1(n1367), .A2(n1368), .A3(n1369), .A4(n1370), .ZN(n1366) );
  NOR4_X1 U801 ( .A1(n1427), .A2(n1428), .A3(n1429), .A4(n1430), .ZN(n1363) );
  NAND4_X1 U802 ( .A1(n1443), .A2(n1444), .A3(n1445), .A4(n1446), .ZN(n1427)
         );
  NAND4_X1 U803 ( .A1(n1439), .A2(n1440), .A3(n1441), .A4(n1442), .ZN(n1428)
         );
  NAND4_X1 U804 ( .A1(n1435), .A2(n1436), .A3(n1437), .A4(n1438), .ZN(n1429)
         );
  INV_X1 U805 ( .I(n1447), .ZN(n580) );
  AOI22_X1 U806 ( .A1(N595), .A2(n484), .B1(n487), .B2(nxt_wr_ptr[63]), .ZN(
        n1447) );
  OAI22_X1 U807 ( .A1(n775), .A2(n457), .B1(n477), .B2(n711), .ZN(n1608) );
  INV_X1 U808 ( .I(N309), .ZN(n711) );
  INV_X1 U809 ( .I(n1272), .ZN(n581) );
  AOI22_X1 U810 ( .A1(N594), .A2(n479), .B1(nxt_wr_ptr[62]), .B2(n489), .ZN(
        n1272) );
  INV_X1 U811 ( .I(n1274), .ZN(n582) );
  AOI22_X1 U812 ( .A1(N593), .A2(n479), .B1(nxt_wr_ptr[61]), .B2(n488), .ZN(
        n1274) );
  INV_X1 U813 ( .I(n1275), .ZN(n583) );
  AOI22_X1 U814 ( .A1(N592), .A2(n479), .B1(nxt_wr_ptr[60]), .B2(n487), .ZN(
        n1275) );
  INV_X1 U815 ( .I(n1276), .ZN(n584) );
  AOI22_X1 U816 ( .A1(N591), .A2(n479), .B1(nxt_wr_ptr[59]), .B2(n486), .ZN(
        n1276) );
  INV_X1 U817 ( .I(n1277), .ZN(n585) );
  AOI22_X1 U818 ( .A1(N590), .A2(n479), .B1(nxt_wr_ptr[58]), .B2(n487), .ZN(
        n1277) );
  INV_X1 U819 ( .I(n1278), .ZN(n586) );
  AOI22_X1 U820 ( .A1(N589), .A2(n479), .B1(nxt_wr_ptr[57]), .B2(n485), .ZN(
        n1278) );
  INV_X1 U821 ( .I(n1279), .ZN(n587) );
  AOI22_X1 U822 ( .A1(N588), .A2(n479), .B1(nxt_wr_ptr[56]), .B2(n487), .ZN(
        n1279) );
  INV_X1 U823 ( .I(n1280), .ZN(n588) );
  AOI22_X1 U824 ( .A1(N587), .A2(n479), .B1(nxt_wr_ptr[55]), .B2(n489), .ZN(
        n1280) );
  INV_X1 U825 ( .I(n1281), .ZN(n589) );
  AOI22_X1 U826 ( .A1(N586), .A2(n479), .B1(nxt_wr_ptr[54]), .B2(n488), .ZN(
        n1281) );
  INV_X1 U827 ( .I(n1282), .ZN(n590) );
  AOI22_X1 U828 ( .A1(N585), .A2(n479), .B1(nxt_wr_ptr[53]), .B2(n485), .ZN(
        n1282) );
  INV_X1 U829 ( .I(n1283), .ZN(n591) );
  AOI22_X1 U830 ( .A1(N584), .A2(n479), .B1(nxt_wr_ptr[52]), .B2(n486), .ZN(
        n1283) );
  INV_X1 U831 ( .I(n1284), .ZN(n592) );
  AOI22_X1 U832 ( .A1(N583), .A2(n479), .B1(nxt_wr_ptr[51]), .B2(n486), .ZN(
        n1284) );
  INV_X1 U833 ( .I(n1285), .ZN(n593) );
  AOI22_X1 U834 ( .A1(N582), .A2(n480), .B1(nxt_wr_ptr[50]), .B2(n486), .ZN(
        n1285) );
  INV_X1 U835 ( .I(n1286), .ZN(n594) );
  AOI22_X1 U836 ( .A1(N581), .A2(n480), .B1(nxt_wr_ptr[49]), .B2(n489), .ZN(
        n1286) );
  INV_X1 U837 ( .I(n1287), .ZN(n595) );
  AOI22_X1 U838 ( .A1(N580), .A2(n480), .B1(nxt_wr_ptr[48]), .B2(n488), .ZN(
        n1287) );
  INV_X1 U839 ( .I(n1288), .ZN(n596) );
  AOI22_X1 U840 ( .A1(N579), .A2(n480), .B1(nxt_wr_ptr[47]), .B2(n486), .ZN(
        n1288) );
  INV_X1 U841 ( .I(n1289), .ZN(n597) );
  AOI22_X1 U842 ( .A1(N578), .A2(n480), .B1(nxt_wr_ptr[46]), .B2(n485), .ZN(
        n1289) );
  INV_X1 U843 ( .I(n1290), .ZN(n598) );
  AOI22_X1 U844 ( .A1(N577), .A2(n480), .B1(nxt_wr_ptr[45]), .B2(n489), .ZN(
        n1290) );
  INV_X1 U845 ( .I(n1291), .ZN(n599) );
  AOI22_X1 U846 ( .A1(N576), .A2(n480), .B1(nxt_wr_ptr[44]), .B2(n488), .ZN(
        n1291) );
  INV_X1 U847 ( .I(n1292), .ZN(n600) );
  AOI22_X1 U848 ( .A1(N575), .A2(n480), .B1(nxt_wr_ptr[43]), .B2(n487), .ZN(
        n1292) );
  INV_X1 U849 ( .I(n1293), .ZN(n601) );
  AOI22_X1 U850 ( .A1(N574), .A2(n480), .B1(nxt_wr_ptr[42]), .B2(n486), .ZN(
        n1293) );
  INV_X1 U851 ( .I(n1294), .ZN(n602) );
  AOI22_X1 U852 ( .A1(N573), .A2(n480), .B1(nxt_wr_ptr[41]), .B2(n485), .ZN(
        n1294) );
  INV_X1 U853 ( .I(n1295), .ZN(n603) );
  AOI22_X1 U854 ( .A1(N572), .A2(n480), .B1(nxt_wr_ptr[40]), .B2(n489), .ZN(
        n1295) );
  INV_X1 U855 ( .I(n1296), .ZN(n604) );
  AOI22_X1 U856 ( .A1(N571), .A2(n480), .B1(nxt_wr_ptr[39]), .B2(n488), .ZN(
        n1296) );
  INV_X1 U857 ( .I(n1297), .ZN(n605) );
  AOI22_X1 U858 ( .A1(N570), .A2(n481), .B1(nxt_wr_ptr[38]), .B2(n485), .ZN(
        n1297) );
  INV_X1 U859 ( .I(n1298), .ZN(n606) );
  AOI22_X1 U860 ( .A1(N569), .A2(n481), .B1(nxt_wr_ptr[37]), .B2(n485), .ZN(
        n1298) );
  INV_X1 U861 ( .I(n1299), .ZN(n607) );
  AOI22_X1 U862 ( .A1(N568), .A2(n481), .B1(nxt_wr_ptr[36]), .B2(n485), .ZN(
        n1299) );
  INV_X1 U863 ( .I(n1300), .ZN(n608) );
  AOI22_X1 U864 ( .A1(N567), .A2(n481), .B1(nxt_wr_ptr[35]), .B2(n485), .ZN(
        n1300) );
  INV_X1 U865 ( .I(n1301), .ZN(n609) );
  AOI22_X1 U866 ( .A1(N566), .A2(n481), .B1(nxt_wr_ptr[34]), .B2(n485), .ZN(
        n1301) );
  INV_X1 U867 ( .I(n1302), .ZN(n610) );
  AOI22_X1 U868 ( .A1(N565), .A2(n481), .B1(nxt_wr_ptr[33]), .B2(n485), .ZN(
        n1302) );
  INV_X1 U869 ( .I(n1303), .ZN(n611) );
  AOI22_X1 U870 ( .A1(N564), .A2(n481), .B1(nxt_wr_ptr[32]), .B2(n485), .ZN(
        n1303) );
  INV_X1 U871 ( .I(n1304), .ZN(n612) );
  AOI22_X1 U872 ( .A1(N563), .A2(n481), .B1(nxt_wr_ptr[31]), .B2(n485), .ZN(
        n1304) );
  INV_X1 U873 ( .I(n1305), .ZN(n613) );
  AOI22_X1 U874 ( .A1(N562), .A2(n481), .B1(nxt_wr_ptr[30]), .B2(n485), .ZN(
        n1305) );
  INV_X1 U875 ( .I(n1306), .ZN(n614) );
  AOI22_X1 U876 ( .A1(N561), .A2(n481), .B1(nxt_wr_ptr[29]), .B2(n485), .ZN(
        n1306) );
  INV_X1 U877 ( .I(n1307), .ZN(n615) );
  AOI22_X1 U878 ( .A1(N560), .A2(n481), .B1(nxt_wr_ptr[28]), .B2(n485), .ZN(
        n1307) );
  INV_X1 U879 ( .I(n1308), .ZN(n616) );
  AOI22_X1 U880 ( .A1(N559), .A2(n481), .B1(nxt_wr_ptr[27]), .B2(n485), .ZN(
        n1308) );
  INV_X1 U881 ( .I(n1309), .ZN(n617) );
  AOI22_X1 U882 ( .A1(N558), .A2(n482), .B1(nxt_wr_ptr[26]), .B2(n486), .ZN(
        n1309) );
  INV_X1 U883 ( .I(n1310), .ZN(n618) );
  AOI22_X1 U884 ( .A1(N557), .A2(n482), .B1(nxt_wr_ptr[25]), .B2(n486), .ZN(
        n1310) );
  INV_X1 U885 ( .I(n1311), .ZN(n619) );
  AOI22_X1 U886 ( .A1(N556), .A2(n482), .B1(nxt_wr_ptr[24]), .B2(n486), .ZN(
        n1311) );
  INV_X1 U887 ( .I(n1312), .ZN(n620) );
  AOI22_X1 U888 ( .A1(N555), .A2(n482), .B1(nxt_wr_ptr[23]), .B2(n486), .ZN(
        n1312) );
  INV_X1 U889 ( .I(n1313), .ZN(n621) );
  AOI22_X1 U890 ( .A1(N554), .A2(n482), .B1(nxt_wr_ptr[22]), .B2(n486), .ZN(
        n1313) );
  INV_X1 U891 ( .I(n1314), .ZN(n622) );
  AOI22_X1 U892 ( .A1(N553), .A2(n482), .B1(nxt_wr_ptr[21]), .B2(n486), .ZN(
        n1314) );
  INV_X1 U893 ( .I(n1315), .ZN(n623) );
  AOI22_X1 U894 ( .A1(N552), .A2(n482), .B1(nxt_wr_ptr[20]), .B2(n486), .ZN(
        n1315) );
  INV_X1 U895 ( .I(n1316), .ZN(n624) );
  AOI22_X1 U896 ( .A1(N551), .A2(n482), .B1(nxt_wr_ptr[19]), .B2(n486), .ZN(
        n1316) );
  INV_X1 U897 ( .I(n1317), .ZN(n625) );
  AOI22_X1 U898 ( .A1(N550), .A2(n482), .B1(nxt_wr_ptr[18]), .B2(n486), .ZN(
        n1317) );
  INV_X1 U899 ( .I(n1318), .ZN(n626) );
  AOI22_X1 U900 ( .A1(N549), .A2(n482), .B1(nxt_wr_ptr[17]), .B2(n486), .ZN(
        n1318) );
  INV_X1 U901 ( .I(n1319), .ZN(n627) );
  AOI22_X1 U902 ( .A1(N548), .A2(n482), .B1(nxt_wr_ptr[16]), .B2(n486), .ZN(
        n1319) );
  NOR2_X1 U903 ( .A1(rst), .A2(n1130), .ZN(n1219) );
  INV_X1 U904 ( .I(n1322), .ZN(n630) );
  AOI22_X1 U905 ( .A1(N545), .A2(n483), .B1(nxt_wr_ptr[13]), .B2(n487), .ZN(
        n1322) );
  INV_X1 U906 ( .I(n1329), .ZN(n637) );
  AOI22_X1 U907 ( .A1(N538), .A2(n483), .B1(nxt_wr_ptr[6]), .B2(n486), .ZN(
        n1329) );
  INV_X1 U908 ( .I(n1321), .ZN(n629) );
  AOI22_X1 U909 ( .A1(N546), .A2(n483), .B1(nxt_wr_ptr[14]), .B2(n489), .ZN(
        n1321) );
  INV_X1 U910 ( .I(n1328), .ZN(n636) );
  AOI22_X1 U911 ( .A1(N539), .A2(n483), .B1(nxt_wr_ptr[7]), .B2(n488), .ZN(
        n1328) );
  INV_X1 U912 ( .I(n1332), .ZN(n640) );
  AOI22_X1 U913 ( .A1(N535), .A2(n483), .B1(nxt_wr_ptr[3]), .B2(n485), .ZN(
        n1332) );
  INV_X1 U914 ( .I(n1320), .ZN(n628) );
  AOI22_X1 U915 ( .A1(N547), .A2(n482), .B1(nxt_wr_ptr[15]), .B2(n486), .ZN(
        n1320) );
  INV_X1 U916 ( .I(n1327), .ZN(n635) );
  AOI22_X1 U917 ( .A1(N540), .A2(n483), .B1(nxt_wr_ptr[8]), .B2(n487), .ZN(
        n1327) );
  INV_X1 U918 ( .I(n1333), .ZN(n641) );
  AOI22_X1 U919 ( .A1(N534), .A2(n484), .B1(nxt_wr_ptr[2]), .B2(n487), .ZN(
        n1333) );
  INV_X1 U920 ( .I(n1326), .ZN(n634) );
  AOI22_X1 U921 ( .A1(N541), .A2(n483), .B1(nxt_wr_ptr[9]), .B2(n486), .ZN(
        n1326) );
  INV_X1 U922 ( .I(n1330), .ZN(n638) );
  AOI22_X1 U923 ( .A1(N537), .A2(n483), .B1(nxt_wr_ptr[5]), .B2(n489), .ZN(
        n1330) );
  INV_X1 U924 ( .I(n1334), .ZN(n642) );
  AOI22_X1 U925 ( .A1(N533), .A2(n484), .B1(nxt_wr_ptr[1]), .B2(n487), .ZN(
        n1334) );
  INV_X1 U926 ( .I(n1323), .ZN(n631) );
  AOI22_X1 U927 ( .A1(N544), .A2(n483), .B1(nxt_wr_ptr[12]), .B2(n488), .ZN(
        n1323) );
  INV_X1 U928 ( .I(n1324), .ZN(n632) );
  AOI22_X1 U929 ( .A1(N543), .A2(n483), .B1(nxt_wr_ptr[11]), .B2(n485), .ZN(
        n1324) );
  INV_X1 U930 ( .I(n1325), .ZN(n633) );
  AOI22_X1 U931 ( .A1(N542), .A2(n483), .B1(nxt_wr_ptr[10]), .B2(n485), .ZN(
        n1325) );
  INV_X1 U932 ( .I(n1331), .ZN(n639) );
  AOI22_X1 U933 ( .A1(N536), .A2(n483), .B1(nxt_wr_ptr[4]), .B2(n487), .ZN(
        n1331) );
  AOI21_X1 U934 ( .A1(n710), .A2(rd), .B(rst), .ZN(n1338) );
  INV_X1 U935 ( .I(rst), .ZN(n1736) );
  NOR2_X1 U936 ( .A1(n571), .A2(rst), .ZN(n978) );
  INV_X1 U937 ( .I(n1012), .ZN(n675) );
  AOI22_X1 U938 ( .A1(N215), .A2(n574), .B1(data_out[33]), .B2(n568), .ZN(
        n1012) );
  INV_X1 U939 ( .I(n1013), .ZN(n674) );
  AOI22_X1 U940 ( .A1(N216), .A2(n574), .B1(data_out[34]), .B2(n568), .ZN(
        n1013) );
  INV_X1 U941 ( .I(n1014), .ZN(n673) );
  AOI22_X1 U942 ( .A1(N217), .A2(n574), .B1(data_out[35]), .B2(n568), .ZN(
        n1014) );
  INV_X1 U943 ( .I(n1011), .ZN(n676) );
  AOI22_X1 U944 ( .A1(N214), .A2(n574), .B1(data_out[32]), .B2(n568), .ZN(
        n1011) );
  INV_X1 U945 ( .I(n1039), .ZN(n648) );
  AOI22_X1 U946 ( .A1(N242), .A2(n577), .B1(data_out[60]), .B2(n571), .ZN(
        n1039) );
  INV_X1 U947 ( .I(n1040), .ZN(n647) );
  AOI22_X1 U948 ( .A1(N243), .A2(n577), .B1(data_out[61]), .B2(n571), .ZN(
        n1040) );
  INV_X1 U949 ( .I(n1041), .ZN(n646) );
  AOI22_X1 U950 ( .A1(N244), .A2(n577), .B1(data_out[62]), .B2(n571), .ZN(
        n1041) );
  INV_X1 U951 ( .I(n1042), .ZN(n645) );
  AOI22_X1 U952 ( .A1(N245), .A2(n577), .B1(data_out[63]), .B2(n571), .ZN(
        n1042) );
  INV_X1 U953 ( .I(n977), .ZN(n708) );
  AOI22_X1 U954 ( .A1(N182), .A2(n572), .B1(data_out[0]), .B2(n566), .ZN(n977)
         );
  INV_X1 U955 ( .I(n980), .ZN(n707) );
  AOI22_X1 U956 ( .A1(N183), .A2(n572), .B1(data_out[1]), .B2(n566), .ZN(n980)
         );
  INV_X1 U957 ( .I(n981), .ZN(n706) );
  AOI22_X1 U958 ( .A1(N184), .A2(n572), .B1(data_out[2]), .B2(n566), .ZN(n981)
         );
  INV_X1 U959 ( .I(n982), .ZN(n705) );
  AOI22_X1 U960 ( .A1(N185), .A2(n572), .B1(data_out[3]), .B2(n566), .ZN(n982)
         );
  INV_X1 U961 ( .I(n983), .ZN(n704) );
  AOI22_X1 U962 ( .A1(N186), .A2(n572), .B1(data_out[4]), .B2(n566), .ZN(n983)
         );
  INV_X1 U963 ( .I(n984), .ZN(n703) );
  AOI22_X1 U964 ( .A1(N187), .A2(n572), .B1(data_out[5]), .B2(n566), .ZN(n984)
         );
  INV_X1 U965 ( .I(n985), .ZN(n702) );
  AOI22_X1 U966 ( .A1(N188), .A2(n572), .B1(data_out[6]), .B2(n566), .ZN(n985)
         );
  INV_X1 U967 ( .I(n986), .ZN(n701) );
  AOI22_X1 U968 ( .A1(N189), .A2(n572), .B1(data_out[7]), .B2(n566), .ZN(n986)
         );
  INV_X1 U969 ( .I(n987), .ZN(n700) );
  AOI22_X1 U970 ( .A1(N190), .A2(n572), .B1(data_out[8]), .B2(n566), .ZN(n987)
         );
  INV_X1 U971 ( .I(n988), .ZN(n699) );
  AOI22_X1 U972 ( .A1(N191), .A2(n572), .B1(data_out[9]), .B2(n566), .ZN(n988)
         );
  INV_X1 U973 ( .I(n989), .ZN(n698) );
  AOI22_X1 U974 ( .A1(N192), .A2(n572), .B1(data_out[10]), .B2(n566), .ZN(n989) );
  INV_X1 U975 ( .I(n990), .ZN(n697) );
  AOI22_X1 U976 ( .A1(N193), .A2(n572), .B1(data_out[11]), .B2(n566), .ZN(n990) );
  INV_X1 U977 ( .I(n991), .ZN(n696) );
  AOI22_X1 U978 ( .A1(N194), .A2(n573), .B1(data_out[12]), .B2(n567), .ZN(n991) );
  INV_X1 U979 ( .I(n992), .ZN(n695) );
  AOI22_X1 U980 ( .A1(N195), .A2(n573), .B1(data_out[13]), .B2(n567), .ZN(n992) );
  INV_X1 U981 ( .I(n993), .ZN(n694) );
  AOI22_X1 U982 ( .A1(N196), .A2(n573), .B1(data_out[14]), .B2(n567), .ZN(n993) );
  INV_X1 U983 ( .I(n994), .ZN(n693) );
  AOI22_X1 U984 ( .A1(N197), .A2(n573), .B1(data_out[15]), .B2(n567), .ZN(n994) );
  INV_X1 U985 ( .I(n995), .ZN(n692) );
  AOI22_X1 U986 ( .A1(N198), .A2(n573), .B1(data_out[16]), .B2(n567), .ZN(n995) );
  INV_X1 U987 ( .I(n996), .ZN(n691) );
  AOI22_X1 U988 ( .A1(N199), .A2(n573), .B1(data_out[17]), .B2(n567), .ZN(n996) );
  INV_X1 U989 ( .I(n997), .ZN(n690) );
  AOI22_X1 U990 ( .A1(N200), .A2(n573), .B1(data_out[18]), .B2(n567), .ZN(n997) );
  INV_X1 U991 ( .I(n998), .ZN(n689) );
  AOI22_X1 U992 ( .A1(N201), .A2(n573), .B1(data_out[19]), .B2(n567), .ZN(n998) );
  INV_X1 U993 ( .I(n999), .ZN(n688) );
  AOI22_X1 U994 ( .A1(N202), .A2(n573), .B1(data_out[20]), .B2(n567), .ZN(n999) );
  INV_X1 U995 ( .I(n1000), .ZN(n687) );
  AOI22_X1 U996 ( .A1(N203), .A2(n573), .B1(data_out[21]), .B2(n567), .ZN(
        n1000) );
  INV_X1 U997 ( .I(n1001), .ZN(n686) );
  AOI22_X1 U998 ( .A1(N204), .A2(n573), .B1(data_out[22]), .B2(n567), .ZN(
        n1001) );
  INV_X1 U999 ( .I(n1002), .ZN(n685) );
  AOI22_X1 U1000 ( .A1(N205), .A2(n573), .B1(data_out[23]), .B2(n567), .ZN(
        n1002) );
  INV_X1 U1001 ( .I(n1003), .ZN(n684) );
  AOI22_X1 U1002 ( .A1(N206), .A2(n574), .B1(data_out[24]), .B2(n568), .ZN(
        n1003) );
  INV_X1 U1003 ( .I(n1004), .ZN(n683) );
  AOI22_X1 U1004 ( .A1(N207), .A2(n574), .B1(data_out[25]), .B2(n568), .ZN(
        n1004) );
  INV_X1 U1005 ( .I(n1005), .ZN(n682) );
  AOI22_X1 U1006 ( .A1(N208), .A2(n574), .B1(data_out[26]), .B2(n568), .ZN(
        n1005) );
  INV_X1 U1007 ( .I(n1006), .ZN(n681) );
  AOI22_X1 U1008 ( .A1(N209), .A2(n574), .B1(data_out[27]), .B2(n568), .ZN(
        n1006) );
  INV_X1 U1009 ( .I(n1007), .ZN(n680) );
  AOI22_X1 U1010 ( .A1(N210), .A2(n574), .B1(data_out[28]), .B2(n568), .ZN(
        n1007) );
  INV_X1 U1011 ( .I(n1008), .ZN(n679) );
  AOI22_X1 U1012 ( .A1(N211), .A2(n574), .B1(data_out[29]), .B2(n568), .ZN(
        n1008) );
  INV_X1 U1013 ( .I(n1009), .ZN(n678) );
  AOI22_X1 U1014 ( .A1(N212), .A2(n574), .B1(data_out[30]), .B2(n568), .ZN(
        n1009) );
  INV_X1 U1015 ( .I(n1010), .ZN(n677) );
  AOI22_X1 U1016 ( .A1(N213), .A2(n574), .B1(data_out[31]), .B2(n568), .ZN(
        n1010) );
  INV_X1 U1017 ( .I(n1020), .ZN(n667) );
  AOI22_X1 U1018 ( .A1(N223), .A2(n575), .B1(data_out[41]), .B2(n569), .ZN(
        n1020) );
  INV_X1 U1019 ( .I(n1015), .ZN(n672) );
  AOI22_X1 U1020 ( .A1(N218), .A2(n575), .B1(data_out[36]), .B2(n569), .ZN(
        n1015) );
  INV_X1 U1021 ( .I(n1017), .ZN(n670) );
  AOI22_X1 U1022 ( .A1(N220), .A2(n575), .B1(data_out[38]), .B2(n569), .ZN(
        n1017) );
  INV_X1 U1023 ( .I(n1021), .ZN(n666) );
  AOI22_X1 U1024 ( .A1(N224), .A2(n575), .B1(data_out[42]), .B2(n569), .ZN(
        n1021) );
  INV_X1 U1025 ( .I(n1023), .ZN(n664) );
  AOI22_X1 U1026 ( .A1(N226), .A2(n575), .B1(data_out[44]), .B2(n569), .ZN(
        n1023) );
  INV_X1 U1027 ( .I(n1025), .ZN(n662) );
  AOI22_X1 U1028 ( .A1(N228), .A2(n575), .B1(data_out[46]), .B2(n569), .ZN(
        n1025) );
  INV_X1 U1029 ( .I(n1018), .ZN(n669) );
  AOI22_X1 U1030 ( .A1(N221), .A2(n575), .B1(data_out[39]), .B2(n569), .ZN(
        n1018) );
  INV_X1 U1031 ( .I(n1026), .ZN(n661) );
  AOI22_X1 U1032 ( .A1(N229), .A2(n575), .B1(data_out[47]), .B2(n569), .ZN(
        n1026) );
  INV_X1 U1033 ( .I(n1016), .ZN(n671) );
  AOI22_X1 U1034 ( .A1(N219), .A2(n575), .B1(data_out[37]), .B2(n569), .ZN(
        n1016) );
  INV_X1 U1035 ( .I(n1022), .ZN(n665) );
  AOI22_X1 U1036 ( .A1(N225), .A2(n575), .B1(data_out[43]), .B2(n569), .ZN(
        n1022) );
  INV_X1 U1037 ( .I(n1024), .ZN(n663) );
  AOI22_X1 U1038 ( .A1(N227), .A2(n575), .B1(data_out[45]), .B2(n569), .ZN(
        n1024) );
  INV_X1 U1039 ( .I(n1019), .ZN(n668) );
  AOI22_X1 U1040 ( .A1(N222), .A2(n575), .B1(data_out[40]), .B2(n569), .ZN(
        n1019) );
  INV_X1 U1041 ( .I(n1027), .ZN(n660) );
  AOI22_X1 U1042 ( .A1(N230), .A2(n576), .B1(data_out[48]), .B2(n570), .ZN(
        n1027) );
  INV_X1 U1043 ( .I(n1028), .ZN(n659) );
  AOI22_X1 U1044 ( .A1(N231), .A2(n576), .B1(data_out[49]), .B2(n570), .ZN(
        n1028) );
  INV_X1 U1045 ( .I(n1029), .ZN(n658) );
  AOI22_X1 U1046 ( .A1(N232), .A2(n576), .B1(data_out[50]), .B2(n570), .ZN(
        n1029) );
  INV_X1 U1047 ( .I(n1030), .ZN(n657) );
  AOI22_X1 U1048 ( .A1(N233), .A2(n576), .B1(data_out[51]), .B2(n570), .ZN(
        n1030) );
  INV_X1 U1049 ( .I(n1031), .ZN(n656) );
  AOI22_X1 U1050 ( .A1(N234), .A2(n576), .B1(data_out[52]), .B2(n570), .ZN(
        n1031) );
  INV_X1 U1051 ( .I(n1032), .ZN(n655) );
  AOI22_X1 U1052 ( .A1(N235), .A2(n576), .B1(data_out[53]), .B2(n570), .ZN(
        n1032) );
  INV_X1 U1053 ( .I(n1033), .ZN(n654) );
  AOI22_X1 U1054 ( .A1(N236), .A2(n576), .B1(data_out[54]), .B2(n570), .ZN(
        n1033) );
  INV_X1 U1055 ( .I(n1034), .ZN(n653) );
  AOI22_X1 U1056 ( .A1(N237), .A2(n576), .B1(data_out[55]), .B2(n570), .ZN(
        n1034) );
  INV_X1 U1057 ( .I(n1035), .ZN(n652) );
  AOI22_X1 U1058 ( .A1(N238), .A2(n576), .B1(data_out[56]), .B2(n570), .ZN(
        n1035) );
  INV_X1 U1059 ( .I(n1036), .ZN(n651) );
  AOI22_X1 U1060 ( .A1(N239), .A2(n576), .B1(data_out[57]), .B2(n570), .ZN(
        n1036) );
  INV_X1 U1061 ( .I(n1037), .ZN(n650) );
  AOI22_X1 U1062 ( .A1(N240), .A2(n576), .B1(data_out[58]), .B2(n570), .ZN(
        n1037) );
  INV_X1 U1063 ( .I(n1038), .ZN(n649) );
  AOI22_X1 U1064 ( .A1(N241), .A2(n576), .B1(data_out[59]), .B2(n570), .ZN(
        n1038) );
  OAI21_X1 U1065 ( .A1(n774), .A2(n478), .B(n1337), .ZN(n1544) );
  NAND2_X1 U1066 ( .A1(rd_ptr[0]), .A2(n1338), .ZN(n1337) );
  INV_X1 U1067 ( .I(n1218), .ZN(n644) );
  AOI22_X1 U1068 ( .A1(n487), .A2(wr_ptr[63]), .B1(n471), .B2(nxt_wr_ptr[63]), 
        .ZN(n1218) );
  INV_X1 U1069 ( .I(n1222), .ZN(n901) );
  AOI22_X1 U1070 ( .A1(n489), .A2(wr_ptr[60]), .B1(n471), .B2(nxt_wr_ptr[60]), 
        .ZN(n1222) );
  INV_X1 U1071 ( .I(n1221), .ZN(n900) );
  AOI22_X1 U1072 ( .A1(n485), .A2(wr_ptr[61]), .B1(n471), .B2(nxt_wr_ptr[61]), 
        .ZN(n1221) );
  INV_X1 U1073 ( .I(n1220), .ZN(n899) );
  AOI22_X1 U1074 ( .A1(n486), .A2(wr_ptr[62]), .B1(n471), .B2(nxt_wr_ptr[62]), 
        .ZN(n1220) );
  INV_X1 U1075 ( .I(full), .ZN(n1712) );
  INV_X1 U1076 ( .I(n1225), .ZN(n904) );
  AOI22_X1 U1077 ( .A1(n486), .A2(wr_ptr[57]), .B1(n470), .B2(nxt_wr_ptr[57]), 
        .ZN(n1225) );
  INV_X1 U1078 ( .I(n1229), .ZN(n908) );
  AOI22_X1 U1079 ( .A1(n489), .A2(wr_ptr[53]), .B1(n470), .B2(nxt_wr_ptr[53]), 
        .ZN(n1229) );
  INV_X1 U1080 ( .I(n1234), .ZN(n912) );
  AOI22_X1 U1081 ( .A1(n489), .A2(wr_ptr[42]), .B1(n470), .B2(nxt_wr_ptr[42]), 
        .ZN(n1234) );
  INV_X1 U1082 ( .I(n1237), .ZN(n915) );
  AOI22_X1 U1083 ( .A1(n489), .A2(wr_ptr[39]), .B1(n469), .B2(nxt_wr_ptr[39]), 
        .ZN(n1237) );
  INV_X1 U1084 ( .I(n1241), .ZN(n919) );
  AOI22_X1 U1085 ( .A1(n489), .A2(wr_ptr[35]), .B1(n469), .B2(nxt_wr_ptr[35]), 
        .ZN(n1241) );
  INV_X1 U1086 ( .I(n1245), .ZN(n923) );
  AOI22_X1 U1087 ( .A1(n488), .A2(wr_ptr[31]), .B1(n469), .B2(nxt_wr_ptr[31]), 
        .ZN(n1245) );
  INV_X1 U1088 ( .I(n1248), .ZN(n926) );
  AOI22_X1 U1089 ( .A1(n488), .A2(wr_ptr[28]), .B1(n468), .B2(nxt_wr_ptr[28]), 
        .ZN(n1248) );
  INV_X1 U1090 ( .I(n1252), .ZN(n930) );
  AOI22_X1 U1091 ( .A1(n488), .A2(wr_ptr[24]), .B1(n468), .B2(nxt_wr_ptr[24]), 
        .ZN(n1252) );
  INV_X1 U1092 ( .I(n1256), .ZN(n934) );
  AOI22_X1 U1093 ( .A1(n488), .A2(wr_ptr[20]), .B1(n468), .B2(nxt_wr_ptr[20]), 
        .ZN(n1256) );
  INV_X1 U1094 ( .I(n1259), .ZN(n937) );
  AOI22_X1 U1095 ( .A1(n488), .A2(wr_ptr[17]), .B1(n468), .B2(nxt_wr_ptr[17]), 
        .ZN(n1259) );
  INV_X1 U1096 ( .I(n1263), .ZN(n941) );
  AOI22_X1 U1097 ( .A1(n487), .A2(wr_ptr[13]), .B1(n467), .B2(nxt_wr_ptr[13]), 
        .ZN(n1263) );
  INV_X1 U1098 ( .I(n1267), .ZN(n945) );
  AOI22_X1 U1099 ( .A1(n487), .A2(wr_ptr[6]), .B1(n467), .B2(nxt_wr_ptr[6]), 
        .ZN(n1267) );
  INV_X1 U1100 ( .I(n1224), .ZN(n903) );
  AOI22_X1 U1101 ( .A1(n489), .A2(wr_ptr[58]), .B1(n470), .B2(nxt_wr_ptr[58]), 
        .ZN(n1224) );
  INV_X1 U1102 ( .I(n1228), .ZN(n907) );
  AOI22_X1 U1103 ( .A1(n489), .A2(wr_ptr[54]), .B1(n470), .B2(nxt_wr_ptr[54]), 
        .ZN(n1228) );
  INV_X1 U1104 ( .I(n1233), .ZN(n911) );
  AOI22_X1 U1105 ( .A1(n489), .A2(wr_ptr[43]), .B1(n470), .B2(nxt_wr_ptr[43]), 
        .ZN(n1233) );
  INV_X1 U1106 ( .I(n1240), .ZN(n918) );
  AOI22_X1 U1107 ( .A1(n489), .A2(wr_ptr[36]), .B1(n469), .B2(nxt_wr_ptr[36]), 
        .ZN(n1240) );
  INV_X1 U1108 ( .I(n1244), .ZN(n922) );
  AOI22_X1 U1109 ( .A1(n489), .A2(wr_ptr[32]), .B1(n469), .B2(nxt_wr_ptr[32]), 
        .ZN(n1244) );
  INV_X1 U1110 ( .I(n1247), .ZN(n925) );
  AOI22_X1 U1111 ( .A1(n488), .A2(wr_ptr[29]), .B1(n469), .B2(nxt_wr_ptr[29]), 
        .ZN(n1247) );
  INV_X1 U1112 ( .I(n1251), .ZN(n929) );
  AOI22_X1 U1113 ( .A1(n488), .A2(wr_ptr[25]), .B1(n468), .B2(nxt_wr_ptr[25]), 
        .ZN(n1251) );
  INV_X1 U1114 ( .I(n1255), .ZN(n933) );
  AOI22_X1 U1115 ( .A1(n488), .A2(wr_ptr[21]), .B1(n468), .B2(nxt_wr_ptr[21]), 
        .ZN(n1255) );
  INV_X1 U1116 ( .I(n1258), .ZN(n936) );
  AOI22_X1 U1117 ( .A1(n488), .A2(wr_ptr[18]), .B1(n468), .B2(nxt_wr_ptr[18]), 
        .ZN(n1258) );
  INV_X1 U1118 ( .I(n1262), .ZN(n940) );
  AOI22_X1 U1119 ( .A1(n487), .A2(wr_ptr[14]), .B1(n467), .B2(nxt_wr_ptr[14]), 
        .ZN(n1262) );
  INV_X1 U1120 ( .I(n1266), .ZN(n944) );
  AOI22_X1 U1121 ( .A1(n487), .A2(wr_ptr[7]), .B1(n467), .B2(nxt_wr_ptr[7]), 
        .ZN(n1266) );
  INV_X1 U1122 ( .I(n1269), .ZN(n947) );
  AOI22_X1 U1123 ( .A1(n487), .A2(wr_ptr[3]), .B1(n467), .B2(nxt_wr_ptr[3]), 
        .ZN(n1269) );
  INV_X1 U1124 ( .I(n1223), .ZN(n902) );
  AOI22_X1 U1125 ( .A1(n488), .A2(wr_ptr[59]), .B1(n470), .B2(nxt_wr_ptr[59]), 
        .ZN(n1223) );
  INV_X1 U1126 ( .I(n1227), .ZN(n906) );
  AOI22_X1 U1127 ( .A1(n485), .A2(wr_ptr[55]), .B1(n470), .B2(nxt_wr_ptr[55]), 
        .ZN(n1227) );
  INV_X1 U1128 ( .I(n1232), .ZN(n910) );
  AOI22_X1 U1129 ( .A1(n489), .A2(wr_ptr[44]), .B1(n470), .B2(nxt_wr_ptr[44]), 
        .ZN(n1232) );
  INV_X1 U1130 ( .I(n1236), .ZN(n914) );
  AOI22_X1 U1131 ( .A1(n489), .A2(wr_ptr[40]), .B1(n469), .B2(nxt_wr_ptr[40]), 
        .ZN(n1236) );
  INV_X1 U1132 ( .I(n1239), .ZN(n917) );
  AOI22_X1 U1133 ( .A1(n489), .A2(wr_ptr[37]), .B1(n469), .B2(nxt_wr_ptr[37]), 
        .ZN(n1239) );
  INV_X1 U1134 ( .I(n1243), .ZN(n921) );
  AOI22_X1 U1135 ( .A1(n489), .A2(wr_ptr[33]), .B1(n469), .B2(nxt_wr_ptr[33]), 
        .ZN(n1243) );
  INV_X1 U1136 ( .I(n1250), .ZN(n928) );
  AOI22_X1 U1137 ( .A1(n488), .A2(wr_ptr[26]), .B1(n468), .B2(nxt_wr_ptr[26]), 
        .ZN(n1250) );
  INV_X1 U1138 ( .I(n1254), .ZN(n932) );
  AOI22_X1 U1139 ( .A1(n488), .A2(wr_ptr[22]), .B1(n468), .B2(nxt_wr_ptr[22]), 
        .ZN(n1254) );
  INV_X1 U1140 ( .I(n1257), .ZN(n935) );
  AOI22_X1 U1141 ( .A1(n488), .A2(wr_ptr[19]), .B1(n468), .B2(nxt_wr_ptr[19]), 
        .ZN(n1257) );
  INV_X1 U1142 ( .I(n1261), .ZN(n939) );
  AOI22_X1 U1143 ( .A1(n488), .A2(wr_ptr[15]), .B1(n467), .B2(nxt_wr_ptr[15]), 
        .ZN(n1261) );
  INV_X1 U1144 ( .I(n1265), .ZN(n943) );
  AOI22_X1 U1145 ( .A1(n487), .A2(wr_ptr[8]), .B1(n467), .B2(nxt_wr_ptr[8]), 
        .ZN(n1265) );
  INV_X1 U1146 ( .I(n1270), .ZN(n948) );
  AOI22_X1 U1147 ( .A1(n487), .A2(wr_ptr[2]), .B1(n467), .B2(nxt_wr_ptr[2]), 
        .ZN(n1270) );
  INV_X1 U1148 ( .I(n1271), .ZN(n949) );
  AOI22_X1 U1149 ( .A1(n487), .A2(wr_ptr[1]), .B1(n467), .B2(nxt_wr_ptr[1]), 
        .ZN(n1271) );
  INV_X1 U1150 ( .I(n1226), .ZN(n905) );
  AOI22_X1 U1151 ( .A1(n485), .A2(wr_ptr[56]), .B1(n470), .B2(nxt_wr_ptr[56]), 
        .ZN(n1226) );
  INV_X1 U1152 ( .I(n1231), .ZN(n909) );
  AOI22_X1 U1153 ( .A1(n489), .A2(wr_ptr[45]), .B1(n470), .B2(nxt_wr_ptr[45]), 
        .ZN(n1231) );
  INV_X1 U1154 ( .I(n1235), .ZN(n913) );
  AOI22_X1 U1155 ( .A1(n489), .A2(wr_ptr[41]), .B1(n470), .B2(nxt_wr_ptr[41]), 
        .ZN(n1235) );
  INV_X1 U1156 ( .I(n1238), .ZN(n916) );
  AOI22_X1 U1157 ( .A1(n489), .A2(wr_ptr[38]), .B1(n469), .B2(nxt_wr_ptr[38]), 
        .ZN(n1238) );
  INV_X1 U1158 ( .I(n1242), .ZN(n920) );
  AOI22_X1 U1159 ( .A1(n489), .A2(wr_ptr[34]), .B1(n469), .B2(nxt_wr_ptr[34]), 
        .ZN(n1242) );
  INV_X1 U1160 ( .I(n1246), .ZN(n924) );
  AOI22_X1 U1161 ( .A1(n488), .A2(wr_ptr[30]), .B1(n469), .B2(nxt_wr_ptr[30]), 
        .ZN(n1246) );
  INV_X1 U1162 ( .I(n1249), .ZN(n927) );
  AOI22_X1 U1163 ( .A1(n488), .A2(wr_ptr[27]), .B1(n468), .B2(nxt_wr_ptr[27]), 
        .ZN(n1249) );
  INV_X1 U1164 ( .I(n1253), .ZN(n931) );
  AOI22_X1 U1165 ( .A1(n488), .A2(wr_ptr[23]), .B1(n468), .B2(nxt_wr_ptr[23]), 
        .ZN(n1253) );
  INV_X1 U1166 ( .I(n1260), .ZN(n938) );
  AOI22_X1 U1167 ( .A1(n488), .A2(wr_ptr[16]), .B1(n467), .B2(nxt_wr_ptr[16]), 
        .ZN(n1260) );
  INV_X1 U1168 ( .I(n1264), .ZN(n942) );
  AOI22_X1 U1169 ( .A1(n487), .A2(wr_ptr[9]), .B1(n467), .B2(nxt_wr_ptr[9]), 
        .ZN(n1264) );
  INV_X1 U1170 ( .I(n1268), .ZN(n946) );
  AOI22_X1 U1171 ( .A1(n487), .A2(wr_ptr[5]), .B1(n467), .B2(nxt_wr_ptr[5]), 
        .ZN(n1268) );
  NAND4_X1 U1172 ( .A1(n1129), .A2(n1130), .A3(wr_ptr[0]), .A4(n1131), .ZN(
        n1065) );
  NOR3_X1 U1173 ( .A1(rst), .A2(wr_ptr[2]), .A3(wr_ptr[1]), .ZN(n1131) );
  INV_X1 U1174 ( .I(n1128), .ZN(n1711) );
  AOI22_X1 U1175 ( .A1(n563), .A2(data_in[0]), .B1(n532), .B2(queue[64]), .ZN(
        n1128) );
  INV_X1 U1176 ( .I(n1127), .ZN(n1710) );
  AOI22_X1 U1177 ( .A1(n563), .A2(data_in[1]), .B1(n532), .B2(queue[65]), .ZN(
        n1127) );
  INV_X1 U1178 ( .I(n1126), .ZN(n1709) );
  AOI22_X1 U1179 ( .A1(n563), .A2(data_in[2]), .B1(n532), .B2(queue[66]), .ZN(
        n1126) );
  INV_X1 U1180 ( .I(n1125), .ZN(n1708) );
  AOI22_X1 U1181 ( .A1(n563), .A2(data_in[3]), .B1(n532), .B2(queue[67]), .ZN(
        n1125) );
  INV_X1 U1182 ( .I(n1124), .ZN(n1707) );
  AOI22_X1 U1183 ( .A1(n562), .A2(data_in[4]), .B1(n532), .B2(queue[68]), .ZN(
        n1124) );
  INV_X1 U1184 ( .I(n1123), .ZN(n1706) );
  AOI22_X1 U1185 ( .A1(n562), .A2(data_in[5]), .B1(n532), .B2(queue[69]), .ZN(
        n1123) );
  INV_X1 U1186 ( .I(n1122), .ZN(n1705) );
  AOI22_X1 U1187 ( .A1(n561), .A2(data_in[6]), .B1(n532), .B2(queue[70]), .ZN(
        n1122) );
  INV_X1 U1188 ( .I(n1121), .ZN(n1704) );
  AOI22_X1 U1189 ( .A1(n561), .A2(data_in[7]), .B1(n532), .B2(queue[71]), .ZN(
        n1121) );
  INV_X1 U1190 ( .I(n1120), .ZN(n1703) );
  AOI22_X1 U1191 ( .A1(n560), .A2(data_in[8]), .B1(n532), .B2(queue[72]), .ZN(
        n1120) );
  INV_X1 U1192 ( .I(n1119), .ZN(n1702) );
  AOI22_X1 U1193 ( .A1(n560), .A2(data_in[9]), .B1(n532), .B2(queue[73]), .ZN(
        n1119) );
  INV_X1 U1194 ( .I(n1118), .ZN(n1701) );
  AOI22_X1 U1195 ( .A1(n559), .A2(data_in[10]), .B1(n532), .B2(queue[74]), 
        .ZN(n1118) );
  INV_X1 U1196 ( .I(n1117), .ZN(n1700) );
  AOI22_X1 U1197 ( .A1(n559), .A2(data_in[11]), .B1(n532), .B2(queue[75]), 
        .ZN(n1117) );
  INV_X1 U1198 ( .I(n1116), .ZN(n1699) );
  AOI22_X1 U1199 ( .A1(n558), .A2(data_in[12]), .B1(n533), .B2(queue[76]), 
        .ZN(n1116) );
  INV_X1 U1200 ( .I(n1115), .ZN(n1698) );
  AOI22_X1 U1201 ( .A1(n558), .A2(data_in[13]), .B1(n533), .B2(queue[77]), 
        .ZN(n1115) );
  INV_X1 U1202 ( .I(n1114), .ZN(n1697) );
  AOI22_X1 U1203 ( .A1(n557), .A2(data_in[14]), .B1(n533), .B2(queue[78]), 
        .ZN(n1114) );
  INV_X1 U1204 ( .I(n1113), .ZN(n1696) );
  AOI22_X1 U1205 ( .A1(n557), .A2(data_in[15]), .B1(n533), .B2(queue[79]), 
        .ZN(n1113) );
  INV_X1 U1206 ( .I(n1112), .ZN(n1695) );
  AOI22_X1 U1207 ( .A1(n556), .A2(data_in[16]), .B1(n533), .B2(queue[80]), 
        .ZN(n1112) );
  INV_X1 U1208 ( .I(n1111), .ZN(n1694) );
  AOI22_X1 U1209 ( .A1(n556), .A2(data_in[17]), .B1(n533), .B2(queue[81]), 
        .ZN(n1111) );
  INV_X1 U1210 ( .I(n1110), .ZN(n1693) );
  AOI22_X1 U1211 ( .A1(n555), .A2(data_in[18]), .B1(n533), .B2(queue[82]), 
        .ZN(n1110) );
  INV_X1 U1212 ( .I(n1109), .ZN(n1692) );
  AOI22_X1 U1213 ( .A1(n555), .A2(data_in[19]), .B1(n533), .B2(queue[83]), 
        .ZN(n1109) );
  INV_X1 U1214 ( .I(n1108), .ZN(n1691) );
  AOI22_X1 U1215 ( .A1(n554), .A2(data_in[20]), .B1(n533), .B2(queue[84]), 
        .ZN(n1108) );
  INV_X1 U1216 ( .I(n1107), .ZN(n1690) );
  AOI22_X1 U1217 ( .A1(n554), .A2(data_in[21]), .B1(n533), .B2(queue[85]), 
        .ZN(n1107) );
  INV_X1 U1218 ( .I(n1106), .ZN(n1689) );
  AOI22_X1 U1219 ( .A1(n553), .A2(data_in[22]), .B1(n533), .B2(queue[86]), 
        .ZN(n1106) );
  INV_X1 U1220 ( .I(n1105), .ZN(n1688) );
  AOI22_X1 U1221 ( .A1(n553), .A2(data_in[23]), .B1(n533), .B2(queue[87]), 
        .ZN(n1105) );
  INV_X1 U1222 ( .I(n1104), .ZN(n1687) );
  AOI22_X1 U1223 ( .A1(n552), .A2(data_in[24]), .B1(n534), .B2(queue[88]), 
        .ZN(n1104) );
  INV_X1 U1224 ( .I(n1103), .ZN(n1686) );
  AOI22_X1 U1225 ( .A1(n552), .A2(data_in[25]), .B1(n534), .B2(queue[89]), 
        .ZN(n1103) );
  INV_X1 U1226 ( .I(n1102), .ZN(n1685) );
  AOI22_X1 U1227 ( .A1(n551), .A2(data_in[26]), .B1(n534), .B2(queue[90]), 
        .ZN(n1102) );
  INV_X1 U1228 ( .I(n1101), .ZN(n1684) );
  AOI22_X1 U1229 ( .A1(n551), .A2(data_in[27]), .B1(n534), .B2(queue[91]), 
        .ZN(n1101) );
  INV_X1 U1230 ( .I(n1100), .ZN(n1683) );
  AOI22_X1 U1231 ( .A1(n550), .A2(data_in[28]), .B1(n534), .B2(queue[92]), 
        .ZN(n1100) );
  INV_X1 U1232 ( .I(n1099), .ZN(n1682) );
  AOI22_X1 U1233 ( .A1(n550), .A2(data_in[29]), .B1(n534), .B2(queue[93]), 
        .ZN(n1099) );
  INV_X1 U1234 ( .I(n1098), .ZN(n1681) );
  AOI22_X1 U1235 ( .A1(n549), .A2(data_in[30]), .B1(n534), .B2(queue[94]), 
        .ZN(n1098) );
  INV_X1 U1236 ( .I(n1097), .ZN(n1680) );
  AOI22_X1 U1237 ( .A1(n549), .A2(data_in[31]), .B1(n534), .B2(queue[95]), 
        .ZN(n1097) );
  INV_X1 U1238 ( .I(n1096), .ZN(n1679) );
  AOI22_X1 U1239 ( .A1(n548), .A2(data_in[32]), .B1(n534), .B2(queue[96]), 
        .ZN(n1096) );
  INV_X1 U1240 ( .I(n1095), .ZN(n1678) );
  AOI22_X1 U1241 ( .A1(n548), .A2(data_in[33]), .B1(n534), .B2(queue[97]), 
        .ZN(n1095) );
  INV_X1 U1242 ( .I(n1094), .ZN(n1677) );
  AOI22_X1 U1243 ( .A1(n547), .A2(data_in[34]), .B1(n534), .B2(queue[98]), 
        .ZN(n1094) );
  INV_X1 U1244 ( .I(n1093), .ZN(n1676) );
  AOI22_X1 U1245 ( .A1(n547), .A2(data_in[35]), .B1(n534), .B2(queue[99]), 
        .ZN(n1093) );
  NAND4_X1 U1246 ( .A1(n1130), .A2(n1736), .A3(n1129), .A4(n1197), .ZN(n1133)
         );
  NOR3_X1 U1247 ( .A1(wr_ptr[0]), .A2(wr_ptr[2]), .A3(wr_ptr[1]), .ZN(n1197)
         );
  INV_X1 U1248 ( .I(n1068), .ZN(n1651) );
  AOI22_X1 U1249 ( .A1(n538), .A2(data_in[60]), .B1(n537), .B2(queue[124]), 
        .ZN(n1068) );
  INV_X1 U1250 ( .I(n1067), .ZN(n1650) );
  AOI22_X1 U1251 ( .A1(n538), .A2(data_in[61]), .B1(n537), .B2(queue[125]), 
        .ZN(n1067) );
  INV_X1 U1252 ( .I(n1066), .ZN(n1649) );
  AOI22_X1 U1253 ( .A1(n538), .A2(data_in[62]), .B1(n537), .B2(queue[126]), 
        .ZN(n1066) );
  INV_X1 U1254 ( .I(n1064), .ZN(n1648) );
  AOI22_X1 U1255 ( .A1(n540), .A2(data_in[63]), .B1(n537), .B2(queue[127]), 
        .ZN(n1064) );
  INV_X1 U1256 ( .I(n1184), .ZN(n1635) );
  AOI22_X1 U1257 ( .A1(data_in[12]), .A2(n524), .B1(n511), .B2(queue[12]), 
        .ZN(n1184) );
  INV_X1 U1258 ( .I(n1183), .ZN(n1634) );
  AOI22_X1 U1259 ( .A1(data_in[13]), .A2(n524), .B1(n510), .B2(queue[13]), 
        .ZN(n1183) );
  INV_X1 U1260 ( .I(n1182), .ZN(n1633) );
  AOI22_X1 U1261 ( .A1(data_in[14]), .A2(n524), .B1(n510), .B2(queue[14]), 
        .ZN(n1182) );
  INV_X1 U1262 ( .I(n1181), .ZN(n1632) );
  AOI22_X1 U1263 ( .A1(data_in[15]), .A2(n524), .B1(n510), .B2(queue[15]), 
        .ZN(n1181) );
  INV_X1 U1264 ( .I(n1180), .ZN(n1631) );
  AOI22_X1 U1265 ( .A1(data_in[16]), .A2(n524), .B1(n509), .B2(queue[16]), 
        .ZN(n1180) );
  INV_X1 U1266 ( .I(n1179), .ZN(n1630) );
  AOI22_X1 U1267 ( .A1(data_in[17]), .A2(n524), .B1(n509), .B2(queue[17]), 
        .ZN(n1179) );
  INV_X1 U1268 ( .I(n1178), .ZN(n1629) );
  AOI22_X1 U1269 ( .A1(data_in[18]), .A2(n524), .B1(n509), .B2(queue[18]), 
        .ZN(n1178) );
  INV_X1 U1270 ( .I(n1177), .ZN(n1628) );
  AOI22_X1 U1271 ( .A1(data_in[19]), .A2(n524), .B1(n508), .B2(queue[19]), 
        .ZN(n1177) );
  INV_X1 U1272 ( .I(n1176), .ZN(n1627) );
  AOI22_X1 U1273 ( .A1(data_in[20]), .A2(n524), .B1(n508), .B2(queue[20]), 
        .ZN(n1176) );
  INV_X1 U1274 ( .I(n1175), .ZN(n1626) );
  AOI22_X1 U1275 ( .A1(data_in[21]), .A2(n524), .B1(n508), .B2(queue[21]), 
        .ZN(n1175) );
  INV_X1 U1276 ( .I(n1174), .ZN(n1625) );
  AOI22_X1 U1277 ( .A1(data_in[22]), .A2(n524), .B1(n507), .B2(queue[22]), 
        .ZN(n1174) );
  INV_X1 U1278 ( .I(n1173), .ZN(n1624) );
  AOI22_X1 U1279 ( .A1(data_in[23]), .A2(n524), .B1(n507), .B2(queue[23]), 
        .ZN(n1173) );
  INV_X1 U1280 ( .I(n1172), .ZN(n1623) );
  AOI22_X1 U1281 ( .A1(data_in[24]), .A2(n524), .B1(n507), .B2(queue[24]), 
        .ZN(n1172) );
  INV_X1 U1282 ( .I(n1171), .ZN(n1622) );
  AOI22_X1 U1283 ( .A1(data_in[25]), .A2(n524), .B1(n506), .B2(queue[25]), 
        .ZN(n1171) );
  INV_X1 U1284 ( .I(n1170), .ZN(n1621) );
  AOI22_X1 U1285 ( .A1(data_in[26]), .A2(n524), .B1(n506), .B2(queue[26]), 
        .ZN(n1170) );
  INV_X1 U1286 ( .I(n1169), .ZN(n1620) );
  AOI22_X1 U1287 ( .A1(data_in[27]), .A2(n524), .B1(n506), .B2(queue[27]), 
        .ZN(n1169) );
  INV_X1 U1288 ( .I(n1168), .ZN(n1619) );
  AOI22_X1 U1289 ( .A1(data_in[28]), .A2(n524), .B1(n505), .B2(queue[28]), 
        .ZN(n1168) );
  INV_X1 U1290 ( .I(n1167), .ZN(n1618) );
  AOI22_X1 U1291 ( .A1(data_in[29]), .A2(n524), .B1(n505), .B2(queue[29]), 
        .ZN(n1167) );
  INV_X1 U1292 ( .I(n1166), .ZN(n1617) );
  AOI22_X1 U1293 ( .A1(data_in[30]), .A2(n524), .B1(n505), .B2(queue[30]), 
        .ZN(n1166) );
  INV_X1 U1294 ( .I(n1165), .ZN(n1616) );
  AOI22_X1 U1295 ( .A1(data_in[31]), .A2(n524), .B1(n504), .B2(queue[31]), 
        .ZN(n1165) );
  INV_X1 U1296 ( .I(n1164), .ZN(n1615) );
  AOI22_X1 U1297 ( .A1(data_in[32]), .A2(n524), .B1(n504), .B2(queue[32]), 
        .ZN(n1164) );
  INV_X1 U1298 ( .I(n1163), .ZN(n1614) );
  AOI22_X1 U1299 ( .A1(data_in[33]), .A2(n524), .B1(n504), .B2(queue[33]), 
        .ZN(n1163) );
  INV_X1 U1300 ( .I(n1162), .ZN(n1613) );
  AOI22_X1 U1301 ( .A1(data_in[34]), .A2(n524), .B1(n503), .B2(queue[34]), 
        .ZN(n1162) );
  INV_X1 U1302 ( .I(n1161), .ZN(n1612) );
  AOI22_X1 U1303 ( .A1(data_in[35]), .A2(n524), .B1(n503), .B2(queue[35]), 
        .ZN(n1161) );
  INV_X1 U1304 ( .I(n1092), .ZN(n1675) );
  AOI22_X1 U1305 ( .A1(n546), .A2(data_in[36]), .B1(n535), .B2(queue[100]), 
        .ZN(n1092) );
  INV_X1 U1306 ( .I(n1091), .ZN(n1674) );
  AOI22_X1 U1307 ( .A1(n546), .A2(data_in[37]), .B1(n535), .B2(queue[101]), 
        .ZN(n1091) );
  INV_X1 U1308 ( .I(n1090), .ZN(n1673) );
  AOI22_X1 U1309 ( .A1(n545), .A2(data_in[38]), .B1(n535), .B2(queue[102]), 
        .ZN(n1090) );
  INV_X1 U1310 ( .I(n1089), .ZN(n1672) );
  AOI22_X1 U1311 ( .A1(n545), .A2(data_in[39]), .B1(n535), .B2(queue[103]), 
        .ZN(n1089) );
  INV_X1 U1312 ( .I(n1088), .ZN(n1671) );
  AOI22_X1 U1313 ( .A1(n544), .A2(data_in[40]), .B1(n535), .B2(queue[104]), 
        .ZN(n1088) );
  INV_X1 U1314 ( .I(n1087), .ZN(n1670) );
  AOI22_X1 U1315 ( .A1(n544), .A2(data_in[41]), .B1(n535), .B2(queue[105]), 
        .ZN(n1087) );
  INV_X1 U1316 ( .I(n1086), .ZN(n1669) );
  AOI22_X1 U1317 ( .A1(n547), .A2(data_in[42]), .B1(n535), .B2(queue[106]), 
        .ZN(n1086) );
  INV_X1 U1318 ( .I(n1085), .ZN(n1668) );
  AOI22_X1 U1319 ( .A1(n546), .A2(data_in[43]), .B1(n535), .B2(queue[107]), 
        .ZN(n1085) );
  INV_X1 U1320 ( .I(n1084), .ZN(n1667) );
  AOI22_X1 U1321 ( .A1(n543), .A2(data_in[44]), .B1(n535), .B2(queue[108]), 
        .ZN(n1084) );
  INV_X1 U1322 ( .I(n1083), .ZN(n1666) );
  AOI22_X1 U1323 ( .A1(n543), .A2(data_in[45]), .B1(n535), .B2(queue[109]), 
        .ZN(n1083) );
  INV_X1 U1324 ( .I(n1082), .ZN(n1665) );
  AOI22_X1 U1325 ( .A1(n542), .A2(data_in[46]), .B1(n535), .B2(queue[110]), 
        .ZN(n1082) );
  INV_X1 U1326 ( .I(n1081), .ZN(n1664) );
  AOI22_X1 U1327 ( .A1(n542), .A2(data_in[47]), .B1(n535), .B2(queue[111]), 
        .ZN(n1081) );
  INV_X1 U1328 ( .I(n1080), .ZN(n1663) );
  AOI22_X1 U1329 ( .A1(n541), .A2(data_in[48]), .B1(n536), .B2(queue[112]), 
        .ZN(n1080) );
  INV_X1 U1330 ( .I(n1079), .ZN(n1662) );
  AOI22_X1 U1331 ( .A1(n541), .A2(data_in[49]), .B1(n536), .B2(queue[113]), 
        .ZN(n1079) );
  INV_X1 U1332 ( .I(n1078), .ZN(n1661) );
  AOI22_X1 U1333 ( .A1(n541), .A2(data_in[50]), .B1(n536), .B2(queue[114]), 
        .ZN(n1078) );
  INV_X1 U1334 ( .I(n1077), .ZN(n1660) );
  AOI22_X1 U1335 ( .A1(n541), .A2(data_in[51]), .B1(n536), .B2(queue[115]), 
        .ZN(n1077) );
  INV_X1 U1336 ( .I(n1076), .ZN(n1659) );
  AOI22_X1 U1337 ( .A1(n543), .A2(data_in[52]), .B1(n536), .B2(queue[116]), 
        .ZN(n1076) );
  INV_X1 U1338 ( .I(n1075), .ZN(n1658) );
  AOI22_X1 U1339 ( .A1(n542), .A2(data_in[53]), .B1(n536), .B2(queue[117]), 
        .ZN(n1075) );
  INV_X1 U1340 ( .I(n1074), .ZN(n1657) );
  AOI22_X1 U1341 ( .A1(n540), .A2(data_in[54]), .B1(n536), .B2(queue[118]), 
        .ZN(n1074) );
  INV_X1 U1342 ( .I(n1073), .ZN(n1656) );
  AOI22_X1 U1343 ( .A1(n540), .A2(data_in[55]), .B1(n536), .B2(queue[119]), 
        .ZN(n1073) );
  INV_X1 U1344 ( .I(n1072), .ZN(n1655) );
  AOI22_X1 U1345 ( .A1(n539), .A2(data_in[56]), .B1(n536), .B2(queue[120]), 
        .ZN(n1072) );
  INV_X1 U1346 ( .I(n1071), .ZN(n1654) );
  AOI22_X1 U1347 ( .A1(n539), .A2(data_in[57]), .B1(n536), .B2(queue[121]), 
        .ZN(n1071) );
  INV_X1 U1348 ( .I(n1070), .ZN(n1653) );
  AOI22_X1 U1349 ( .A1(n539), .A2(data_in[58]), .B1(n536), .B2(queue[122]), 
        .ZN(n1070) );
  INV_X1 U1350 ( .I(n1069), .ZN(n1652) );
  AOI22_X1 U1351 ( .A1(n538), .A2(data_in[59]), .B1(n536), .B2(queue[123]), 
        .ZN(n1069) );
  INV_X1 U1352 ( .I(n1196), .ZN(n1647) );
  AOI22_X1 U1353 ( .A1(data_in[0]), .A2(n524), .B1(n515), .B2(queue[0]), .ZN(
        n1196) );
  INV_X1 U1354 ( .I(n1136), .ZN(n954) );
  AOI22_X1 U1355 ( .A1(data_in[60]), .A2(n524), .B1(n495), .B2(queue[60]), 
        .ZN(n1136) );
  INV_X1 U1356 ( .I(n1135), .ZN(n953) );
  AOI22_X1 U1357 ( .A1(data_in[61]), .A2(n524), .B1(n494), .B2(queue[61]), 
        .ZN(n1135) );
  INV_X1 U1358 ( .I(n1134), .ZN(n952) );
  AOI22_X1 U1359 ( .A1(data_in[62]), .A2(n524), .B1(n494), .B2(queue[62]), 
        .ZN(n1134) );
  INV_X1 U1360 ( .I(n1132), .ZN(n951) );
  AOI22_X1 U1361 ( .A1(data_in[63]), .A2(n524), .B1(n494), .B2(queue[63]), 
        .ZN(n1132) );
  INV_X1 U1362 ( .I(n1195), .ZN(n1646) );
  AOI22_X1 U1363 ( .A1(data_in[1]), .A2(n524), .B1(n514), .B2(queue[1]), .ZN(
        n1195) );
  INV_X1 U1364 ( .I(n1194), .ZN(n1645) );
  AOI22_X1 U1365 ( .A1(data_in[2]), .A2(n524), .B1(n514), .B2(queue[2]), .ZN(
        n1194) );
  INV_X1 U1366 ( .I(n1193), .ZN(n1644) );
  AOI22_X1 U1367 ( .A1(data_in[3]), .A2(n524), .B1(n514), .B2(queue[3]), .ZN(
        n1193) );
  INV_X1 U1368 ( .I(n1192), .ZN(n1643) );
  AOI22_X1 U1369 ( .A1(data_in[4]), .A2(n524), .B1(n513), .B2(queue[4]), .ZN(
        n1192) );
  INV_X1 U1370 ( .I(n1191), .ZN(n1642) );
  AOI22_X1 U1371 ( .A1(data_in[5]), .A2(n524), .B1(n513), .B2(queue[5]), .ZN(
        n1191) );
  INV_X1 U1372 ( .I(n1190), .ZN(n1641) );
  AOI22_X1 U1373 ( .A1(data_in[6]), .A2(n524), .B1(n513), .B2(queue[6]), .ZN(
        n1190) );
  INV_X1 U1374 ( .I(n1189), .ZN(n1640) );
  AOI22_X1 U1375 ( .A1(data_in[7]), .A2(n524), .B1(n512), .B2(queue[7]), .ZN(
        n1189) );
  INV_X1 U1376 ( .I(n1188), .ZN(n1639) );
  AOI22_X1 U1377 ( .A1(data_in[8]), .A2(n524), .B1(n512), .B2(queue[8]), .ZN(
        n1188) );
  INV_X1 U1378 ( .I(n1187), .ZN(n1638) );
  AOI22_X1 U1379 ( .A1(data_in[9]), .A2(n524), .B1(n512), .B2(queue[9]), .ZN(
        n1187) );
  INV_X1 U1380 ( .I(n1186), .ZN(n1637) );
  AOI22_X1 U1381 ( .A1(data_in[10]), .A2(n524), .B1(n511), .B2(queue[10]), 
        .ZN(n1186) );
  INV_X1 U1382 ( .I(n1185), .ZN(n1636) );
  AOI22_X1 U1383 ( .A1(data_in[11]), .A2(n524), .B1(n511), .B2(queue[11]), 
        .ZN(n1185) );
  INV_X1 U1384 ( .I(n1160), .ZN(n1611) );
  AOI22_X1 U1385 ( .A1(data_in[36]), .A2(n524), .B1(n503), .B2(queue[36]), 
        .ZN(n1160) );
  INV_X1 U1386 ( .I(n1159), .ZN(n1336) );
  AOI22_X1 U1387 ( .A1(data_in[37]), .A2(n524), .B1(n502), .B2(queue[37]), 
        .ZN(n1159) );
  INV_X1 U1388 ( .I(n1158), .ZN(n976) );
  AOI22_X1 U1389 ( .A1(data_in[38]), .A2(n524), .B1(n502), .B2(queue[38]), 
        .ZN(n1158) );
  INV_X1 U1390 ( .I(n1157), .ZN(n975) );
  AOI22_X1 U1391 ( .A1(data_in[39]), .A2(n524), .B1(n502), .B2(queue[39]), 
        .ZN(n1157) );
  INV_X1 U1392 ( .I(n1156), .ZN(n974) );
  AOI22_X1 U1393 ( .A1(data_in[40]), .A2(n524), .B1(n501), .B2(queue[40]), 
        .ZN(n1156) );
  INV_X1 U1394 ( .I(n1155), .ZN(n973) );
  AOI22_X1 U1395 ( .A1(data_in[41]), .A2(n524), .B1(n501), .B2(queue[41]), 
        .ZN(n1155) );
  INV_X1 U1396 ( .I(n1154), .ZN(n972) );
  AOI22_X1 U1397 ( .A1(data_in[42]), .A2(n524), .B1(n501), .B2(queue[42]), 
        .ZN(n1154) );
  INV_X1 U1398 ( .I(n1153), .ZN(n971) );
  AOI22_X1 U1399 ( .A1(data_in[43]), .A2(n524), .B1(n500), .B2(queue[43]), 
        .ZN(n1153) );
  INV_X1 U1400 ( .I(n1152), .ZN(n970) );
  AOI22_X1 U1401 ( .A1(data_in[44]), .A2(n524), .B1(n500), .B2(queue[44]), 
        .ZN(n1152) );
  INV_X1 U1402 ( .I(n1151), .ZN(n969) );
  AOI22_X1 U1403 ( .A1(data_in[45]), .A2(n524), .B1(n500), .B2(queue[45]), 
        .ZN(n1151) );
  INV_X1 U1404 ( .I(n1150), .ZN(n968) );
  AOI22_X1 U1405 ( .A1(data_in[46]), .A2(n524), .B1(n499), .B2(queue[46]), 
        .ZN(n1150) );
  INV_X1 U1406 ( .I(n1149), .ZN(n967) );
  AOI22_X1 U1407 ( .A1(data_in[47]), .A2(n524), .B1(n499), .B2(queue[47]), 
        .ZN(n1149) );
  INV_X1 U1408 ( .I(n1148), .ZN(n966) );
  AOI22_X1 U1409 ( .A1(data_in[48]), .A2(n524), .B1(n499), .B2(queue[48]), 
        .ZN(n1148) );
  INV_X1 U1410 ( .I(n1147), .ZN(n965) );
  AOI22_X1 U1411 ( .A1(data_in[49]), .A2(n524), .B1(n498), .B2(queue[49]), 
        .ZN(n1147) );
  INV_X1 U1412 ( .I(n1146), .ZN(n964) );
  AOI22_X1 U1413 ( .A1(data_in[50]), .A2(n524), .B1(n498), .B2(queue[50]), 
        .ZN(n1146) );
  INV_X1 U1414 ( .I(n1145), .ZN(n963) );
  AOI22_X1 U1415 ( .A1(data_in[51]), .A2(n524), .B1(n498), .B2(queue[51]), 
        .ZN(n1145) );
  INV_X1 U1416 ( .I(n1144), .ZN(n962) );
  AOI22_X1 U1417 ( .A1(data_in[52]), .A2(n524), .B1(n497), .B2(queue[52]), 
        .ZN(n1144) );
  INV_X1 U1418 ( .I(n1143), .ZN(n961) );
  AOI22_X1 U1419 ( .A1(data_in[53]), .A2(n524), .B1(n497), .B2(queue[53]), 
        .ZN(n1143) );
  INV_X1 U1420 ( .I(n1142), .ZN(n960) );
  AOI22_X1 U1421 ( .A1(data_in[54]), .A2(n524), .B1(n497), .B2(queue[54]), 
        .ZN(n1142) );
  INV_X1 U1422 ( .I(n1141), .ZN(n959) );
  AOI22_X1 U1423 ( .A1(data_in[55]), .A2(n524), .B1(n496), .B2(queue[55]), 
        .ZN(n1141) );
  INV_X1 U1424 ( .I(n1140), .ZN(n958) );
  AOI22_X1 U1425 ( .A1(data_in[56]), .A2(n524), .B1(n496), .B2(queue[56]), 
        .ZN(n1140) );
  INV_X1 U1426 ( .I(n1139), .ZN(n957) );
  AOI22_X1 U1427 ( .A1(data_in[57]), .A2(n524), .B1(n496), .B2(queue[57]), 
        .ZN(n1139) );
  INV_X1 U1428 ( .I(n1138), .ZN(n956) );
  AOI22_X1 U1429 ( .A1(data_in[58]), .A2(n524), .B1(n495), .B2(queue[58]), 
        .ZN(n1138) );
  INV_X1 U1430 ( .I(n1137), .ZN(n955) );
  AOI22_X1 U1431 ( .A1(data_in[59]), .A2(n524), .B1(n495), .B2(queue[59]), 
        .ZN(n1137) );
  INV_X1 U1432 ( .I(empty), .ZN(n710) );
  OAI22_X1 U1433 ( .A1(n491), .A2(n643), .B1(n487), .B2(n1449), .ZN(n1610) );
  AOI21_X1 U1434 ( .A1(N532), .A2(n1448), .B(rst), .ZN(n1449) );
  INV_X1 U1435 ( .I(rd_ptr[56]), .ZN(n885) );
  OAI22_X1 U1436 ( .A1(n774), .A2(n457), .B1(n1338), .B2(n1340), .ZN(n1607) );
  AOI21_X1 U1437 ( .A1(N246), .A2(n1341), .B(rst), .ZN(n1340) );
  NOR4_X1 U1438 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1198)
         );
  NOR4_X1 U1439 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199)
         );
  INV_X1 U1440 ( .I(rd_ptr[5]), .ZN(n783) );
  INV_X1 U1441 ( .I(rd_ptr[63]), .ZN(n898) );
  INV_X1 U1442 ( .I(rd_ptr[41]), .ZN(n855) );
  INV_X1 U1443 ( .I(rd_ptr[45]), .ZN(n863) );
  INV_X1 U1444 ( .I(rd_ptr[49]), .ZN(n871) );
  INV_X1 U1445 ( .I(rd_ptr[26]), .ZN(n825) );
  INV_X1 U1446 ( .I(rd_ptr[30]), .ZN(n833) );
  INV_X1 U1447 ( .I(rd_ptr[54]), .ZN(n881) );
  INV_X1 U1448 ( .I(rd_ptr[58]), .ZN(n889) );
  INV_X1 U1449 ( .I(rd_ptr[3]), .ZN(n779) );
  INV_X1 U1450 ( .I(rd_ptr[55]), .ZN(n883) );
  INV_X1 U1451 ( .I(rd_ptr[59]), .ZN(n891) );
  INV_X1 U1452 ( .I(rd_ptr[62]), .ZN(n897) );
  INV_X1 U1453 ( .I(rd_ptr[40]), .ZN(n853) );
  INV_X1 U1454 ( .I(rd_ptr[44]), .ZN(n861) );
  INV_X1 U1455 ( .I(rd_ptr[25]), .ZN(n823) );
  INV_X1 U1456 ( .I(rd_ptr[29]), .ZN(n831) );
  OAI22_X1 U1457 ( .A1(n1713), .A2(n490), .B1(n456), .B2(n643), .ZN(n1481) );
  INV_X1 U1458 ( .I(wr_ptr[0]), .ZN(n1713) );
  INV_X1 U1459 ( .I(rd_ptr[53]), .ZN(n879) );
  INV_X1 U1460 ( .I(rd_ptr[57]), .ZN(n887) );
  INV_X1 U1461 ( .I(rd_ptr[39]), .ZN(n851) );
  INV_X1 U1462 ( .I(rd_ptr[42]), .ZN(n857) );
  INV_X1 U1463 ( .I(rd_ptr[9]), .ZN(n791) );
  INV_X1 U1464 ( .I(rd_ptr[52]), .ZN(n877) );
  INV_X1 U1465 ( .I(rd_ptr[34]), .ZN(n841) );
  INV_X1 U1466 ( .I(rd_ptr[38]), .ZN(n849) );
  INV_X1 U1467 ( .I(rd_ptr[14]), .ZN(n801) );
  INV_X1 U1468 ( .I(rd_ptr[18]), .ZN(n809) );
  INV_X1 U1469 ( .I(rd_ptr[61]), .ZN(n895) );
  INV_X1 U1470 ( .I(rd_ptr[43]), .ZN(n859) );
  INV_X1 U1471 ( .I(rd_ptr[47]), .ZN(n867) );
  INV_X1 U1472 ( .I(rd_ptr[24]), .ZN(n821) );
  INV_X1 U1473 ( .I(rd_ptr[28]), .ZN(n829) );
  INV_X1 U1474 ( .I(rd_ptr[32]), .ZN(n837) );
  INV_X1 U1475 ( .I(rd_ptr[8]), .ZN(n789) );
  INV_X1 U1476 ( .I(rd_ptr[48]), .ZN(n869) );
  INV_X1 U1477 ( .I(rd_ptr[51]), .ZN(n875) );
  INV_X1 U1478 ( .I(rd_ptr[33]), .ZN(n839) );
  INV_X1 U1479 ( .I(rd_ptr[13]), .ZN(n799) );
  INV_X1 U1480 ( .I(rd_ptr[17]), .ZN(n807) );
  NAND3_X1 U1481 ( .A1(n710), .A2(n793), .A3(rd), .ZN(n1063) );
  INV_X1 U1482 ( .I(rd_ptr[60]), .ZN(n893) );
  INV_X1 U1483 ( .I(rd_ptr[6]), .ZN(n785) );
  INV_X1 U1484 ( .I(rd_ptr[46]), .ZN(n865) );
  INV_X1 U1485 ( .I(rd_ptr[23]), .ZN(n819) );
  INV_X1 U1486 ( .I(rd_ptr[27]), .ZN(n827) );
  INV_X1 U1487 ( .I(rd_ptr[31]), .ZN(n835) );
  INV_X1 U1488 ( .I(rd_ptr[11]), .ZN(n795) );
  INV_X1 U1489 ( .I(rd_ptr[22]), .ZN(n817) );
  INV_X1 U1490 ( .I(rd_ptr[7]), .ZN(n787) );
  INV_X1 U1491 ( .I(rd_ptr[50]), .ZN(n873) );
  INV_X1 U1492 ( .I(rd_ptr[36]), .ZN(n845) );
  INV_X1 U1493 ( .I(rd_ptr[12]), .ZN(n797) );
  INV_X1 U1494 ( .I(rd_ptr[16]), .ZN(n805) );
  INV_X1 U1495 ( .I(rd_ptr[37]), .ZN(n847) );
  INV_X1 U1496 ( .I(rd_ptr[21]), .ZN(n815) );
  INV_X1 U1497 ( .I(rd_ptr[10]), .ZN(n793) );
  INV_X1 U1498 ( .I(rd_ptr[4]), .ZN(n781) );
  INV_X1 U1499 ( .I(rd_ptr[35]), .ZN(n843) );
  INV_X1 U1500 ( .I(rd_ptr[15]), .ZN(n803) );
  INV_X1 U1501 ( .I(rd_ptr[20]), .ZN(n813) );
  NAND4_X1 U1502 ( .A1(n1719), .A2(n1721), .A3(n1717), .A4(n1213), .ZN(n1210)
         );
  NOR4_X1 U1503 ( .A1(wr_ptr[16]), .A2(wr_ptr[15]), .A3(wr_ptr[14]), .A4(
        wr_ptr[13]), .ZN(n1213) );
  INV_X1 U1504 ( .I(rd_ptr[19]), .ZN(n811) );
  NOR4_X1 U1505 ( .A1(wr_ptr[9]), .A2(wr_ptr[8]), .A3(wr_ptr[7]), .A4(
        wr_ptr[6]), .ZN(n1208) );
  NOR4_X1 U1506 ( .A1(wr_ptr[39]), .A2(wr_ptr[38]), .A3(wr_ptr[37]), .A4(
        wr_ptr[36]), .ZN(n1217) );
  NAND4_X1 U1507 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1200)
         );
  NOR4_X1 U1508 ( .A1(wr_ptr[56]), .A2(wr_ptr[55]), .A3(wr_ptr[54]), .A4(
        wr_ptr[53]), .ZN(n1205) );
  NOR4_X1 U1509 ( .A1(wr_ptr[5]), .A2(wr_ptr[59]), .A3(wr_ptr[58]), .A4(
        wr_ptr[57]), .ZN(n1206) );
  NOR4_X1 U1510 ( .A1(wr_ptr[63]), .A2(wr_ptr[62]), .A3(wr_ptr[61]), .A4(
        wr_ptr[60]), .ZN(n1207) );
  NAND4_X1 U1511 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1209)
         );
  NOR3_X1 U1512 ( .A1(wr_ptr[25]), .A2(wr_ptr[27]), .A3(wr_ptr[26]), .ZN(n1214) );
  NOR4_X1 U1513 ( .A1(wr_ptr[31]), .A2(wr_ptr[30]), .A3(wr_ptr[29]), .A4(
        wr_ptr[28]), .ZN(n1215) );
  NOR4_X1 U1514 ( .A1(wr_ptr[35]), .A2(wr_ptr[34]), .A3(wr_ptr[33]), .A4(
        wr_ptr[32]), .ZN(n1216) );
  INV_X1 U1515 ( .I(wr_ptr[49]), .ZN(n1729) );
  INV_X1 U1516 ( .I(wr_ptr[52]), .ZN(n1735) );
  INV_X1 U1517 ( .I(wr_ptr[47]), .ZN(n1725) );
  INV_X1 U1518 ( .I(wr_ptr[50]), .ZN(n1731) );
  INV_X1 U1519 ( .I(wr_ptr[48]), .ZN(n1727) );
  INV_X1 U1520 ( .I(wr_ptr[51]), .ZN(n1733) );
  INV_X1 U1521 ( .I(wr_ptr[10]), .ZN(n1717) );
  INV_X1 U1522 ( .I(wr_ptr[46]), .ZN(n1723) );
  INV_X1 U1523 ( .I(wr_ptr[4]), .ZN(n1715) );
  INV_X1 U1524 ( .I(wr_ptr[12]), .ZN(n1721) );
  INV_X1 U1525 ( .I(wr_ptr[11]), .ZN(n1719) );
  NOR4_X1 U1526 ( .A1(n1454), .A2(n1455), .A3(n1456), .A4(n1457), .ZN(n1453)
         );
  NAND4_X1 U1527 ( .A1(nxt_wr_ptr[0]), .A2(n1716), .A3(n1718), .A4(n1720), 
        .ZN(n1469) );
  INV_X1 U1614 ( .I(nxt_wr_ptr[49]), .ZN(n1728) );
  INV_X1 U1615 ( .I(nxt_wr_ptr[12]), .ZN(n1720) );
  INV_X1 U1616 ( .I(nxt_wr_ptr[48]), .ZN(n1726) );
  INV_X1 U1617 ( .I(nxt_wr_ptr[11]), .ZN(n1718) );
  INV_X1 U1618 ( .I(nxt_wr_ptr[46]), .ZN(n1722) );
  INV_X1 U1619 ( .I(nxt_wr_ptr[47]), .ZN(n1724) );
  INV_X1 U1620 ( .I(nxt_wr_ptr[50]), .ZN(n1730) );
  INV_X1 U1621 ( .I(nxt_wr_ptr[10]), .ZN(n1716) );
  INV_X1 U1622 ( .I(nxt_wr_ptr[52]), .ZN(n1734) );
  INV_X1 U1623 ( .I(nxt_wr_ptr[51]), .ZN(n1732) );
  INV_X1 U1624 ( .I(nxt_wr_ptr[4]), .ZN(n1714) );
  INV_X1 U1625 ( .I(nxt_rd_ptr[63]), .ZN(n775) );
  INV_X1 U1626 ( .I(nxt_rd_ptr[5]), .ZN(n782) );
  INV_X1 U1627 ( .I(nxt_rd_ptr[56]), .ZN(n884) );
  INV_X1 U1628 ( .I(nxt_rd_ptr[41]), .ZN(n854) );
  INV_X1 U1629 ( .I(nxt_rd_ptr[55]), .ZN(n882) );
  NAND4_X1 U1630 ( .A1(nxt_rd_ptr[0]), .A2(n792), .A3(n794), .A4(n796), .ZN(
        n1361) );
  INV_X1 U1631 ( .I(nxt_rd_ptr[27]), .ZN(n826) );
  INV_X1 U1632 ( .I(nxt_rd_ptr[12]), .ZN(n796) );
  INV_X1 U1633 ( .I(nxt_rd_ptr[49]), .ZN(n870) );
  INV_X1 U1634 ( .I(nxt_rd_ptr[34]), .ZN(n840) );
  INV_X1 U1635 ( .I(nxt_rd_ptr[45]), .ZN(n862) );
  INV_X1 U1636 ( .I(nxt_rd_ptr[30]), .ZN(n832) );
  INV_X1 U1637 ( .I(nxt_rd_ptr[11]), .ZN(n794) );
  INV_X1 U1638 ( .I(nxt_rd_ptr[48]), .ZN(n868) );
  INV_X1 U1639 ( .I(nxt_rd_ptr[62]), .ZN(n896) );
  INV_X1 U1640 ( .I(nxt_rd_ptr[59]), .ZN(n890) );
  INV_X1 U1641 ( .I(nxt_rd_ptr[33]), .ZN(n838) );
  INV_X1 U1642 ( .I(nxt_rd_ptr[40]), .ZN(n852) );
  INV_X1 U1643 ( .I(nxt_rd_ptr[44]), .ZN(n860) );
  INV_X1 U1644 ( .I(nxt_rd_ptr[26]), .ZN(n824) );
  INV_X1 U1645 ( .I(nxt_rd_ptr[43]), .ZN(n858) );
  INV_X1 U1646 ( .I(nxt_rd_ptr[3]), .ZN(n778) );
  INV_X1 U1647 ( .I(nxt_rd_ptr[54]), .ZN(n880) );
  INV_X1 U1648 ( .I(nxt_rd_ptr[61]), .ZN(n894) );
  INV_X1 U1649 ( .I(nxt_rd_ptr[58]), .ZN(n888) );
  INV_X1 U1650 ( .I(nxt_rd_ptr[25]), .ZN(n822) );
  INV_X1 U1651 ( .I(nxt_rd_ptr[29]), .ZN(n830) );
  INV_X1 U1652 ( .I(nxt_rd_ptr[53]), .ZN(n878) );
  INV_X1 U1653 ( .I(nxt_rd_ptr[9]), .ZN(n790) );
  INV_X1 U1654 ( .I(nxt_rd_ptr[52]), .ZN(n876) );
  INV_X1 U1655 ( .I(nxt_rd_ptr[38]), .ZN(n848) );
  INV_X1 U1656 ( .I(nxt_rd_ptr[16]), .ZN(n804) );
  INV_X1 U1657 ( .I(nxt_rd_ptr[51]), .ZN(n874) );
  INV_X1 U1658 ( .I(nxt_rd_ptr[15]), .ZN(n802) );
  INV_X1 U1659 ( .I(nxt_rd_ptr[19]), .ZN(n810) );
  INV_X1 U1660 ( .I(nxt_rd_ptr[8]), .ZN(n788) );
  INV_X1 U1661 ( .I(nxt_rd_ptr[37]), .ZN(n846) );
  INV_X1 U1662 ( .I(nxt_rd_ptr[47]), .ZN(n866) );
  INV_X1 U1663 ( .I(nxt_rd_ptr[10]), .ZN(n792) );
  INV_X1 U1664 ( .I(nxt_rd_ptr[14]), .ZN(n800) );
  INV_X1 U1665 ( .I(nxt_rd_ptr[7]), .ZN(n786) );
  INV_X1 U1666 ( .I(nxt_rd_ptr[50]), .ZN(n872) );
  INV_X1 U1667 ( .I(nxt_rd_ptr[32]), .ZN(n836) );
  INV_X1 U1668 ( .I(nxt_rd_ptr[18]), .ZN(n808) );
  INV_X1 U1669 ( .I(nxt_rd_ptr[39]), .ZN(n850) );
  INV_X1 U1670 ( .I(nxt_rd_ptr[31]), .ZN(n834) );
  INV_X1 U1671 ( .I(nxt_rd_ptr[60]), .ZN(n892) );
  INV_X1 U1672 ( .I(nxt_rd_ptr[57]), .ZN(n886) );
  INV_X1 U1673 ( .I(nxt_rd_ptr[42]), .ZN(n856) );
  INV_X1 U1674 ( .I(nxt_rd_ptr[46]), .ZN(n864) );
  INV_X1 U1675 ( .I(nxt_rd_ptr[24]), .ZN(n820) );
  INV_X1 U1676 ( .I(nxt_rd_ptr[28]), .ZN(n828) );
  INV_X1 U1677 ( .I(nxt_rd_ptr[2]), .ZN(n777) );
  INV_X1 U1678 ( .I(nxt_rd_ptr[23]), .ZN(n818) );
  INV_X1 U1679 ( .I(nxt_rd_ptr[22]), .ZN(n816) );
  INV_X1 U1680 ( .I(nxt_rd_ptr[36]), .ZN(n844) );
  INV_X1 U1681 ( .I(nxt_rd_ptr[21]), .ZN(n814) );
  INV_X1 U1682 ( .I(nxt_rd_ptr[4]), .ZN(n780) );
  INV_X1 U1683 ( .I(nxt_rd_ptr[35]), .ZN(n842) );
  INV_X1 U1684 ( .I(nxt_rd_ptr[13]), .ZN(n798) );
  INV_X1 U1685 ( .I(nxt_rd_ptr[6]), .ZN(n784) );
  INV_X1 U1686 ( .I(nxt_rd_ptr[17]), .ZN(n806) );
  INV_X1 U1687 ( .I(nxt_rd_ptr[1]), .ZN(n776) );
  INV_X1 U1688 ( .I(nxt_rd_ptr[20]), .ZN(n812) );
  NAND4_X1 U1689 ( .A1(n1431), .A2(n1432), .A3(n1433), .A4(n1434), .ZN(n1430)
         );
  INV_X1 U1690 ( .I(nxt_rd_ptr[0]), .ZN(n774) );
  NAND4_X1 U1691 ( .A1(n1411), .A2(n1412), .A3(n1413), .A4(n1414), .ZN(n1410)
         );
  NAND4_X1 U1692 ( .A1(n1391), .A2(n1392), .A3(n1393), .A4(n1394), .ZN(n1390)
         );
  NAND4_X1 U1693 ( .A1(n1371), .A2(n1372), .A3(n1373), .A4(n1374), .ZN(n1370)
         );
  NAND4_X1 U1694 ( .A1(n1395), .A2(n1396), .A3(n1397), .A4(n1398), .ZN(n1389)
         );
  NAND4_X1 U1695 ( .A1(n1375), .A2(n1376), .A3(n1377), .A4(n1378), .ZN(n1369)
         );
  NAND4_X1 U1696 ( .A1(n1383), .A2(n1384), .A3(n1385), .A4(n1386), .ZN(n1367)
         );
  NAND4_X1 U1697 ( .A1(n1415), .A2(n1416), .A3(n1417), .A4(n1418), .ZN(n1409)
         );
  NAND4_X1 U1698 ( .A1(n1379), .A2(n1380), .A3(n1381), .A4(n1382), .ZN(n1368)
         );
  NAND4_X1 U1699 ( .A1(n1399), .A2(n1400), .A3(n1401), .A4(n1402), .ZN(n1388)
         );
  NAND4_X1 U1700 ( .A1(n1419), .A2(n1420), .A3(n1421), .A4(n1422), .ZN(n1408)
         );
  BUF_X2 U1701 ( .I(rd_ptr[0]), .Z(n450) );
  NAND4_X1 U1702 ( .A1(n1403), .A2(n1404), .A3(n1405), .A4(n1406), .ZN(n1387)
         );
  NAND4_X1 U1703 ( .A1(n1423), .A2(n1424), .A3(n1425), .A4(n1426), .ZN(n1407)
         );
  BUF_X2 U1704 ( .I(rd_ptr[0]), .Z(n455) );
  BUF_X2 U1705 ( .I(rd_ptr[0]), .Z(n454) );
  BUF_X2 U1706 ( .I(rd_ptr[0]), .Z(n453) );
  BUF_X2 U1707 ( .I(rd_ptr[0]), .Z(n452) );
  BUF_X2 U1708 ( .I(rd_ptr[0]), .Z(n451) );
  INV_X1 U1709 ( .I(nxt_wr_ptr[0]), .ZN(n643) );
  MUX2_X1 U1710 ( .I0(queue[0]), .I1(queue[64]), .S(n455), .Z(N182) );
  MUX2_X1 U1711 ( .I0(queue[1]), .I1(queue[65]), .S(n455), .Z(N183) );
  MUX2_X1 U1712 ( .I0(queue[2]), .I1(queue[66]), .S(n455), .Z(N184) );
  MUX2_X1 U1713 ( .I0(queue[3]), .I1(queue[67]), .S(n455), .Z(N185) );
  MUX2_X1 U1714 ( .I0(queue[4]), .I1(queue[68]), .S(n455), .Z(N186) );
  MUX2_X1 U1715 ( .I0(queue[5]), .I1(queue[69]), .S(n455), .Z(N187) );
  MUX2_X1 U1716 ( .I0(queue[6]), .I1(queue[70]), .S(n455), .Z(N188) );
  MUX2_X1 U1717 ( .I0(queue[7]), .I1(queue[71]), .S(n455), .Z(N189) );
  MUX2_X1 U1718 ( .I0(queue[8]), .I1(queue[72]), .S(n455), .Z(N190) );
  MUX2_X1 U1719 ( .I0(queue[9]), .I1(queue[73]), .S(n455), .Z(N191) );
  MUX2_X1 U1720 ( .I0(queue[10]), .I1(queue[74]), .S(n455), .Z(N192) );
  MUX2_X1 U1721 ( .I0(queue[11]), .I1(queue[75]), .S(n455), .Z(N193) );
  MUX2_X1 U1722 ( .I0(queue[12]), .I1(queue[76]), .S(n454), .Z(N194) );
  MUX2_X1 U1723 ( .I0(queue[13]), .I1(queue[77]), .S(n454), .Z(N195) );
  MUX2_X1 U1724 ( .I0(queue[14]), .I1(queue[78]), .S(n454), .Z(N196) );
  MUX2_X1 U1725 ( .I0(queue[15]), .I1(queue[79]), .S(n454), .Z(N197) );
  MUX2_X1 U1726 ( .I0(queue[16]), .I1(queue[80]), .S(n454), .Z(N198) );
  MUX2_X1 U1727 ( .I0(queue[17]), .I1(queue[81]), .S(n454), .Z(N199) );
  MUX2_X1 U1728 ( .I0(queue[18]), .I1(queue[82]), .S(n454), .Z(N200) );
  MUX2_X1 U1729 ( .I0(queue[19]), .I1(queue[83]), .S(n454), .Z(N201) );
  MUX2_X1 U1730 ( .I0(queue[20]), .I1(queue[84]), .S(n454), .Z(N202) );
  MUX2_X1 U1731 ( .I0(queue[21]), .I1(queue[85]), .S(n454), .Z(N203) );
  MUX2_X1 U1732 ( .I0(queue[22]), .I1(queue[86]), .S(n454), .Z(N204) );
  MUX2_X1 U1733 ( .I0(queue[23]), .I1(queue[87]), .S(n454), .Z(N205) );
  MUX2_X1 U1734 ( .I0(queue[24]), .I1(queue[88]), .S(n453), .Z(N206) );
  MUX2_X1 U1735 ( .I0(queue[25]), .I1(queue[89]), .S(n453), .Z(N207) );
  MUX2_X1 U1736 ( .I0(queue[26]), .I1(queue[90]), .S(n453), .Z(N208) );
  MUX2_X1 U1737 ( .I0(queue[27]), .I1(queue[91]), .S(n453), .Z(N209) );
  MUX2_X1 U1738 ( .I0(queue[28]), .I1(queue[92]), .S(n453), .Z(N210) );
  MUX2_X1 U1739 ( .I0(queue[29]), .I1(queue[93]), .S(n453), .Z(N211) );
  MUX2_X1 U1740 ( .I0(queue[30]), .I1(queue[94]), .S(n453), .Z(N212) );
  MUX2_X1 U1741 ( .I0(queue[31]), .I1(queue[95]), .S(n453), .Z(N213) );
  MUX2_X1 U1742 ( .I0(queue[32]), .I1(queue[96]), .S(n453), .Z(N214) );
  MUX2_X1 U1743 ( .I0(queue[33]), .I1(queue[97]), .S(n453), .Z(N215) );
  MUX2_X1 U1744 ( .I0(queue[34]), .I1(queue[98]), .S(n453), .Z(N216) );
  MUX2_X1 U1745 ( .I0(queue[35]), .I1(queue[99]), .S(n453), .Z(N217) );
  MUX2_X1 U1746 ( .I0(queue[36]), .I1(queue[100]), .S(n452), .Z(N218) );
  MUX2_X1 U1747 ( .I0(queue[37]), .I1(queue[101]), .S(n452), .Z(N219) );
  MUX2_X1 U1748 ( .I0(queue[38]), .I1(queue[102]), .S(n452), .Z(N220) );
  MUX2_X1 U1749 ( .I0(queue[39]), .I1(queue[103]), .S(n452), .Z(N221) );
  MUX2_X1 U1750 ( .I0(queue[40]), .I1(queue[104]), .S(n452), .Z(N222) );
  MUX2_X1 U1751 ( .I0(queue[41]), .I1(queue[105]), .S(n452), .Z(N223) );
  MUX2_X1 U1752 ( .I0(queue[42]), .I1(queue[106]), .S(n452), .Z(N224) );
  MUX2_X1 U1753 ( .I0(queue[43]), .I1(queue[107]), .S(n452), .Z(N225) );
  MUX2_X1 U1754 ( .I0(queue[44]), .I1(queue[108]), .S(n452), .Z(N226) );
  MUX2_X1 U1755 ( .I0(queue[45]), .I1(queue[109]), .S(n452), .Z(N227) );
  MUX2_X1 U1756 ( .I0(queue[46]), .I1(queue[110]), .S(n452), .Z(N228) );
  MUX2_X1 U1757 ( .I0(queue[47]), .I1(queue[111]), .S(n452), .Z(N229) );
  MUX2_X1 U1758 ( .I0(queue[48]), .I1(queue[112]), .S(n451), .Z(N230) );
  MUX2_X1 U1759 ( .I0(queue[49]), .I1(queue[113]), .S(n451), .Z(N231) );
  MUX2_X1 U1760 ( .I0(queue[50]), .I1(queue[114]), .S(n451), .Z(N232) );
  MUX2_X1 U1761 ( .I0(queue[51]), .I1(queue[115]), .S(n451), .Z(N233) );
  MUX2_X1 U1762 ( .I0(queue[52]), .I1(queue[116]), .S(n451), .Z(N234) );
  MUX2_X1 U1763 ( .I0(queue[53]), .I1(queue[117]), .S(n451), .Z(N235) );
  MUX2_X1 U1764 ( .I0(queue[54]), .I1(queue[118]), .S(n451), .Z(N236) );
  MUX2_X1 U1765 ( .I0(queue[55]), .I1(queue[119]), .S(n451), .Z(N237) );
  MUX2_X1 U1766 ( .I0(queue[56]), .I1(queue[120]), .S(n451), .Z(N238) );
  MUX2_X1 U1767 ( .I0(queue[57]), .I1(queue[121]), .S(n451), .Z(N239) );
  MUX2_X1 U1768 ( .I0(queue[58]), .I1(queue[122]), .S(n451), .Z(N240) );
  MUX2_X1 U1769 ( .I0(queue[59]), .I1(queue[123]), .S(n451), .Z(N241) );
  MUX2_X1 U1770 ( .I0(queue[60]), .I1(queue[124]), .S(n450), .Z(N242) );
  MUX2_X1 U1771 ( .I0(queue[61]), .I1(queue[125]), .S(n450), .Z(N243) );
  MUX2_X1 U1772 ( .I0(queue[62]), .I1(queue[126]), .S(n450), .Z(N244) );
  MUX2_X1 U1773 ( .I0(queue[63]), .I1(queue[127]), .S(n450), .Z(N245) );
  INV_X1 U1774 ( .I(n565), .ZN(n537) );
  INV_X1 U1775 ( .I(n525), .ZN(n538) );
  INV_X1 U1776 ( .I(n525), .ZN(n539) );
  INV_X1 U1777 ( .I(n525), .ZN(n540) );
  INV_X1 U1778 ( .I(n526), .ZN(n541) );
  INV_X1 U1779 ( .I(n526), .ZN(n542) );
  INV_X1 U1780 ( .I(n526), .ZN(n543) );
  INV_X1 U1781 ( .I(n527), .ZN(n544) );
  INV_X1 U1782 ( .I(n527), .ZN(n545) );
  INV_X1 U1783 ( .I(n527), .ZN(n546) );
  INV_X1 U1784 ( .I(n527), .ZN(n547) );
  INV_X1 U1785 ( .I(n528), .ZN(n548) );
  INV_X1 U1786 ( .I(n528), .ZN(n549) );
  INV_X1 U1787 ( .I(n528), .ZN(n550) );
  INV_X1 U1788 ( .I(n528), .ZN(n551) );
  INV_X1 U1789 ( .I(n528), .ZN(n552) );
  INV_X1 U1790 ( .I(n529), .ZN(n553) );
  INV_X1 U1791 ( .I(n529), .ZN(n554) );
  INV_X1 U1792 ( .I(n529), .ZN(n555) );
  INV_X1 U1793 ( .I(n529), .ZN(n556) );
  INV_X1 U1794 ( .I(n529), .ZN(n557) );
  INV_X1 U1795 ( .I(n530), .ZN(n558) );
  INV_X1 U1796 ( .I(n530), .ZN(n559) );
  INV_X1 U1797 ( .I(n530), .ZN(n560) );
  INV_X1 U1798 ( .I(n530), .ZN(n561) );
  INV_X1 U1799 ( .I(n530), .ZN(n562) );
  INV_X1 U1800 ( .I(n531), .ZN(n563) );
  INV_X1 U1801 ( .I(n531), .ZN(n564) );
  INV_X1 U1802 ( .I(n531), .ZN(n565) );
endmodule


module circ_q_WORD_SZ64_0_DW01_inc_0 ( A, SUM );
  input [63:0] A;
  output [63:0] SUM;

  wire   [63:2] carry;

  HA_X1 U1_1_62 ( .A(A[62]), .B(carry[62]), .CO(carry[63]), .S(SUM[62]) );
  HA_X1 U1_1_61 ( .A(A[61]), .B(carry[61]), .CO(carry[62]), .S(SUM[61]) );
  HA_X1 U1_1_60 ( .A(A[60]), .B(carry[60]), .CO(carry[61]), .S(SUM[60]) );
  HA_X1 U1_1_59 ( .A(A[59]), .B(carry[59]), .CO(carry[60]), .S(SUM[59]) );
  HA_X1 U1_1_58 ( .A(A[58]), .B(carry[58]), .CO(carry[59]), .S(SUM[58]) );
  HA_X1 U1_1_57 ( .A(A[57]), .B(carry[57]), .CO(carry[58]), .S(SUM[57]) );
  HA_X1 U1_1_56 ( .A(A[56]), .B(carry[56]), .CO(carry[57]), .S(SUM[56]) );
  HA_X1 U1_1_55 ( .A(A[55]), .B(carry[55]), .CO(carry[56]), .S(SUM[55]) );
  HA_X1 U1_1_54 ( .A(A[54]), .B(carry[54]), .CO(carry[55]), .S(SUM[54]) );
  HA_X1 U1_1_53 ( .A(A[53]), .B(carry[53]), .CO(carry[54]), .S(SUM[53]) );
  HA_X1 U1_1_52 ( .A(A[52]), .B(carry[52]), .CO(carry[53]), .S(SUM[52]) );
  HA_X1 U1_1_51 ( .A(A[51]), .B(carry[51]), .CO(carry[52]), .S(SUM[51]) );
  HA_X1 U1_1_50 ( .A(A[50]), .B(carry[50]), .CO(carry[51]), .S(SUM[50]) );
  HA_X1 U1_1_49 ( .A(A[49]), .B(carry[49]), .CO(carry[50]), .S(SUM[49]) );
  HA_X1 U1_1_48 ( .A(A[48]), .B(carry[48]), .CO(carry[49]), .S(SUM[48]) );
  HA_X1 U1_1_47 ( .A(A[47]), .B(carry[47]), .CO(carry[48]), .S(SUM[47]) );
  HA_X1 U1_1_46 ( .A(A[46]), .B(carry[46]), .CO(carry[47]), .S(SUM[46]) );
  HA_X1 U1_1_45 ( .A(A[45]), .B(carry[45]), .CO(carry[46]), .S(SUM[45]) );
  HA_X1 U1_1_44 ( .A(A[44]), .B(carry[44]), .CO(carry[45]), .S(SUM[44]) );
  HA_X1 U1_1_43 ( .A(A[43]), .B(carry[43]), .CO(carry[44]), .S(SUM[43]) );
  HA_X1 U1_1_42 ( .A(A[42]), .B(carry[42]), .CO(carry[43]), .S(SUM[42]) );
  HA_X1 U1_1_41 ( .A(A[41]), .B(carry[41]), .CO(carry[42]), .S(SUM[41]) );
  HA_X1 U1_1_40 ( .A(A[40]), .B(carry[40]), .CO(carry[41]), .S(SUM[40]) );
  HA_X1 U1_1_39 ( .A(A[39]), .B(carry[39]), .CO(carry[40]), .S(SUM[39]) );
  HA_X1 U1_1_38 ( .A(A[38]), .B(carry[38]), .CO(carry[39]), .S(SUM[38]) );
  HA_X1 U1_1_37 ( .A(A[37]), .B(carry[37]), .CO(carry[38]), .S(SUM[37]) );
  HA_X1 U1_1_36 ( .A(A[36]), .B(carry[36]), .CO(carry[37]), .S(SUM[36]) );
  HA_X1 U1_1_35 ( .A(A[35]), .B(carry[35]), .CO(carry[36]), .S(SUM[35]) );
  HA_X1 U1_1_34 ( .A(A[34]), .B(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  HA_X1 U1_1_33 ( .A(A[33]), .B(carry[33]), .CO(carry[34]), .S(SUM[33]) );
  HA_X1 U1_1_32 ( .A(A[32]), .B(carry[32]), .CO(carry[33]), .S(SUM[32]) );
  HA_X1 U1_1_31 ( .A(A[31]), .B(carry[31]), .CO(carry[32]), .S(SUM[31]) );
  HA_X1 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A1(carry[63]), .A2(A[63]), .Z(SUM[63]) );
endmodule


module circ_q_WORD_SZ64_0_DW01_inc_1 ( A, SUM );
  input [63:0] A;
  output [63:0] SUM;

  wire   [63:2] carry;

  HA_X1 U1_1_62 ( .A(A[62]), .B(carry[62]), .CO(carry[63]), .S(SUM[62]) );
  HA_X1 U1_1_61 ( .A(A[61]), .B(carry[61]), .CO(carry[62]), .S(SUM[61]) );
  HA_X1 U1_1_60 ( .A(A[60]), .B(carry[60]), .CO(carry[61]), .S(SUM[60]) );
  HA_X1 U1_1_59 ( .A(A[59]), .B(carry[59]), .CO(carry[60]), .S(SUM[59]) );
  HA_X1 U1_1_58 ( .A(A[58]), .B(carry[58]), .CO(carry[59]), .S(SUM[58]) );
  HA_X1 U1_1_57 ( .A(A[57]), .B(carry[57]), .CO(carry[58]), .S(SUM[57]) );
  HA_X1 U1_1_56 ( .A(A[56]), .B(carry[56]), .CO(carry[57]), .S(SUM[56]) );
  HA_X1 U1_1_55 ( .A(A[55]), .B(carry[55]), .CO(carry[56]), .S(SUM[55]) );
  HA_X1 U1_1_54 ( .A(A[54]), .B(carry[54]), .CO(carry[55]), .S(SUM[54]) );
  HA_X1 U1_1_53 ( .A(A[53]), .B(carry[53]), .CO(carry[54]), .S(SUM[53]) );
  HA_X1 U1_1_52 ( .A(A[52]), .B(carry[52]), .CO(carry[53]), .S(SUM[52]) );
  HA_X1 U1_1_51 ( .A(A[51]), .B(carry[51]), .CO(carry[52]), .S(SUM[51]) );
  HA_X1 U1_1_50 ( .A(A[50]), .B(carry[50]), .CO(carry[51]), .S(SUM[50]) );
  HA_X1 U1_1_49 ( .A(A[49]), .B(carry[49]), .CO(carry[50]), .S(SUM[49]) );
  HA_X1 U1_1_48 ( .A(A[48]), .B(carry[48]), .CO(carry[49]), .S(SUM[48]) );
  HA_X1 U1_1_47 ( .A(A[47]), .B(carry[47]), .CO(carry[48]), .S(SUM[47]) );
  HA_X1 U1_1_46 ( .A(A[46]), .B(carry[46]), .CO(carry[47]), .S(SUM[46]) );
  HA_X1 U1_1_45 ( .A(A[45]), .B(carry[45]), .CO(carry[46]), .S(SUM[45]) );
  HA_X1 U1_1_44 ( .A(A[44]), .B(carry[44]), .CO(carry[45]), .S(SUM[44]) );
  HA_X1 U1_1_43 ( .A(A[43]), .B(carry[43]), .CO(carry[44]), .S(SUM[43]) );
  HA_X1 U1_1_42 ( .A(A[42]), .B(carry[42]), .CO(carry[43]), .S(SUM[42]) );
  HA_X1 U1_1_41 ( .A(A[41]), .B(carry[41]), .CO(carry[42]), .S(SUM[41]) );
  HA_X1 U1_1_40 ( .A(A[40]), .B(carry[40]), .CO(carry[41]), .S(SUM[40]) );
  HA_X1 U1_1_39 ( .A(A[39]), .B(carry[39]), .CO(carry[40]), .S(SUM[39]) );
  HA_X1 U1_1_38 ( .A(A[38]), .B(carry[38]), .CO(carry[39]), .S(SUM[38]) );
  HA_X1 U1_1_37 ( .A(A[37]), .B(carry[37]), .CO(carry[38]), .S(SUM[37]) );
  HA_X1 U1_1_36 ( .A(A[36]), .B(carry[36]), .CO(carry[37]), .S(SUM[36]) );
  HA_X1 U1_1_35 ( .A(A[35]), .B(carry[35]), .CO(carry[36]), .S(SUM[35]) );
  HA_X1 U1_1_34 ( .A(A[34]), .B(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  HA_X1 U1_1_33 ( .A(A[33]), .B(carry[33]), .CO(carry[34]), .S(SUM[33]) );
  HA_X1 U1_1_32 ( .A(A[32]), .B(carry[32]), .CO(carry[33]), .S(SUM[32]) );
  HA_X1 U1_1_31 ( .A(A[31]), .B(carry[31]), .CO(carry[32]), .S(SUM[31]) );
  HA_X1 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A1(carry[63]), .A2(A[63]), .Z(SUM[63]) );
endmodule


module circ_q_WORD_SZ64_0 ( clk, rst, rd, wr, full, empty, data_in, data_out
 );
  input [63:0] data_in;
  output [63:0] data_out;
  input clk, rst, rd, wr;
  output full, empty;
  wire   N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192,
         N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280,
         N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291,
         N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302,
         N303, N304, N305, N306, N307, N308, N309, N532, N533, N534, N535,
         N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546,
         N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557,
         N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568,
         N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579,
         N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590,
         N591, N592, N593, N594, N595, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n1336, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369;
  wire   [63:0] nxt_wr_ptr;
  wire   [63:0] nxt_rd_ptr;
  wire   [63:0] rd_ptr;
  wire   [63:0] wr_ptr;
  wire   [127:0] queue;

  DFFSNQ_X1 nxt_wr_ptr_reg_0_ ( .D(n1737), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[0]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_63_ ( .D(n580), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[63]) );
  DFFSNQ_X1 empty_reg ( .D(n1738), .CLK(clk), .SN(1'b1), .Q(empty) );
  DFFSNQ_X1 nxt_rd_ptr_reg_0_ ( .D(n1740), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[0]) );
  DFFSNQ_X1 rd_ptr_reg_0_ ( .D(n1803), .CLK(clk), .SN(1'b1), .Q(rd_ptr[0]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_63_ ( .D(n1739), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[63]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_1_ ( .D(n1741), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[1]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_2_ ( .D(n1742), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[2]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_3_ ( .D(n1743), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[3]) );
  DFFSNQ_X1 rd_ptr_reg_3_ ( .D(n1804), .CLK(clk), .SN(1'b1), .Q(rd_ptr[3]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_4_ ( .D(n1744), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[4]) );
  DFFSNQ_X1 rd_ptr_reg_4_ ( .D(n1805), .CLK(clk), .SN(1'b1), .Q(rd_ptr[4]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_5_ ( .D(n1745), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[5]) );
  DFFSNQ_X1 rd_ptr_reg_5_ ( .D(n1806), .CLK(clk), .SN(1'b1), .Q(rd_ptr[5]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_6_ ( .D(n1746), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[6]) );
  DFFSNQ_X1 rd_ptr_reg_6_ ( .D(n1807), .CLK(clk), .SN(1'b1), .Q(rd_ptr[6]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_7_ ( .D(n1747), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[7]) );
  DFFSNQ_X1 rd_ptr_reg_7_ ( .D(n1808), .CLK(clk), .SN(1'b1), .Q(rd_ptr[7]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_8_ ( .D(n1748), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[8]) );
  DFFSNQ_X1 rd_ptr_reg_8_ ( .D(n1809), .CLK(clk), .SN(1'b1), .Q(rd_ptr[8]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_9_ ( .D(n1749), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[9]) );
  DFFSNQ_X1 rd_ptr_reg_9_ ( .D(n1810), .CLK(clk), .SN(1'b1), .Q(rd_ptr[9]) );
  DFFSNQ_X1 nxt_rd_ptr_reg_10_ ( .D(n1750), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[10]) );
  DFFSNQ_X1 rd_ptr_reg_10_ ( .D(n1811), .CLK(clk), .SN(1'b1), .Q(rd_ptr[10])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_11_ ( .D(n1751), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[11]) );
  DFFSNQ_X1 rd_ptr_reg_11_ ( .D(n1812), .CLK(clk), .SN(1'b1), .Q(rd_ptr[11])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_12_ ( .D(n1752), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[12]) );
  DFFSNQ_X1 rd_ptr_reg_12_ ( .D(n1813), .CLK(clk), .SN(1'b1), .Q(rd_ptr[12])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_13_ ( .D(n1753), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[13]) );
  DFFSNQ_X1 rd_ptr_reg_13_ ( .D(n1814), .CLK(clk), .SN(1'b1), .Q(rd_ptr[13])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_14_ ( .D(n1754), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[14]) );
  DFFSNQ_X1 rd_ptr_reg_14_ ( .D(n1815), .CLK(clk), .SN(1'b1), .Q(rd_ptr[14])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_15_ ( .D(n1755), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[15]) );
  DFFSNQ_X1 rd_ptr_reg_15_ ( .D(n1816), .CLK(clk), .SN(1'b1), .Q(rd_ptr[15])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_16_ ( .D(n1756), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[16]) );
  DFFSNQ_X1 rd_ptr_reg_16_ ( .D(n1817), .CLK(clk), .SN(1'b1), .Q(rd_ptr[16])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_17_ ( .D(n1757), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[17]) );
  DFFSNQ_X1 rd_ptr_reg_17_ ( .D(n1818), .CLK(clk), .SN(1'b1), .Q(rd_ptr[17])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_18_ ( .D(n1758), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[18]) );
  DFFSNQ_X1 rd_ptr_reg_18_ ( .D(n1819), .CLK(clk), .SN(1'b1), .Q(rd_ptr[18])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_19_ ( .D(n1759), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[19]) );
  DFFSNQ_X1 rd_ptr_reg_19_ ( .D(n1820), .CLK(clk), .SN(1'b1), .Q(rd_ptr[19])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_20_ ( .D(n1760), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[20]) );
  DFFSNQ_X1 rd_ptr_reg_20_ ( .D(n1821), .CLK(clk), .SN(1'b1), .Q(rd_ptr[20])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_21_ ( .D(n1761), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[21]) );
  DFFSNQ_X1 rd_ptr_reg_21_ ( .D(n1822), .CLK(clk), .SN(1'b1), .Q(rd_ptr[21])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_22_ ( .D(n1762), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[22]) );
  DFFSNQ_X1 rd_ptr_reg_22_ ( .D(n1823), .CLK(clk), .SN(1'b1), .Q(rd_ptr[22])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_23_ ( .D(n1763), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[23]) );
  DFFSNQ_X1 rd_ptr_reg_23_ ( .D(n1824), .CLK(clk), .SN(1'b1), .Q(rd_ptr[23])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_24_ ( .D(n1764), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[24]) );
  DFFSNQ_X1 rd_ptr_reg_24_ ( .D(n1825), .CLK(clk), .SN(1'b1), .Q(rd_ptr[24])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_25_ ( .D(n1765), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[25]) );
  DFFSNQ_X1 rd_ptr_reg_25_ ( .D(n1826), .CLK(clk), .SN(1'b1), .Q(rd_ptr[25])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_26_ ( .D(n1766), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[26]) );
  DFFSNQ_X1 rd_ptr_reg_26_ ( .D(n1827), .CLK(clk), .SN(1'b1), .Q(rd_ptr[26])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_27_ ( .D(n1767), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[27]) );
  DFFSNQ_X1 rd_ptr_reg_27_ ( .D(n1828), .CLK(clk), .SN(1'b1), .Q(rd_ptr[27])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_28_ ( .D(n1768), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[28]) );
  DFFSNQ_X1 rd_ptr_reg_28_ ( .D(n1829), .CLK(clk), .SN(1'b1), .Q(rd_ptr[28])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_29_ ( .D(n1769), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[29]) );
  DFFSNQ_X1 rd_ptr_reg_29_ ( .D(n1830), .CLK(clk), .SN(1'b1), .Q(rd_ptr[29])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_30_ ( .D(n1770), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[30]) );
  DFFSNQ_X1 rd_ptr_reg_30_ ( .D(n1831), .CLK(clk), .SN(1'b1), .Q(rd_ptr[30])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_31_ ( .D(n1771), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[31]) );
  DFFSNQ_X1 rd_ptr_reg_31_ ( .D(n1832), .CLK(clk), .SN(1'b1), .Q(rd_ptr[31])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_32_ ( .D(n1772), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[32]) );
  DFFSNQ_X1 rd_ptr_reg_32_ ( .D(n1833), .CLK(clk), .SN(1'b1), .Q(rd_ptr[32])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_33_ ( .D(n1773), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[33]) );
  DFFSNQ_X1 rd_ptr_reg_33_ ( .D(n1834), .CLK(clk), .SN(1'b1), .Q(rd_ptr[33])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_34_ ( .D(n1774), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[34]) );
  DFFSNQ_X1 rd_ptr_reg_34_ ( .D(n1835), .CLK(clk), .SN(1'b1), .Q(rd_ptr[34])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_35_ ( .D(n1775), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[35]) );
  DFFSNQ_X1 rd_ptr_reg_35_ ( .D(n1836), .CLK(clk), .SN(1'b1), .Q(rd_ptr[35])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_36_ ( .D(n1776), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[36]) );
  DFFSNQ_X1 rd_ptr_reg_36_ ( .D(n1837), .CLK(clk), .SN(1'b1), .Q(rd_ptr[36])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_37_ ( .D(n1777), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[37]) );
  DFFSNQ_X1 rd_ptr_reg_37_ ( .D(n1838), .CLK(clk), .SN(1'b1), .Q(rd_ptr[37])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_38_ ( .D(n1778), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[38]) );
  DFFSNQ_X1 rd_ptr_reg_38_ ( .D(n1839), .CLK(clk), .SN(1'b1), .Q(rd_ptr[38])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_39_ ( .D(n1779), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[39]) );
  DFFSNQ_X1 rd_ptr_reg_39_ ( .D(n1840), .CLK(clk), .SN(1'b1), .Q(rd_ptr[39])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_40_ ( .D(n1780), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[40]) );
  DFFSNQ_X1 rd_ptr_reg_40_ ( .D(n1841), .CLK(clk), .SN(1'b1), .Q(rd_ptr[40])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_41_ ( .D(n1781), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[41]) );
  DFFSNQ_X1 rd_ptr_reg_41_ ( .D(n1842), .CLK(clk), .SN(1'b1), .Q(rd_ptr[41])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_42_ ( .D(n1782), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[42]) );
  DFFSNQ_X1 rd_ptr_reg_42_ ( .D(n1843), .CLK(clk), .SN(1'b1), .Q(rd_ptr[42])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_43_ ( .D(n1783), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[43]) );
  DFFSNQ_X1 rd_ptr_reg_43_ ( .D(n1844), .CLK(clk), .SN(1'b1), .Q(rd_ptr[43])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_44_ ( .D(n1784), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[44]) );
  DFFSNQ_X1 rd_ptr_reg_44_ ( .D(n1845), .CLK(clk), .SN(1'b1), .Q(rd_ptr[44])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_45_ ( .D(n1785), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[45]) );
  DFFSNQ_X1 rd_ptr_reg_45_ ( .D(n1846), .CLK(clk), .SN(1'b1), .Q(rd_ptr[45])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_46_ ( .D(n1786), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[46]) );
  DFFSNQ_X1 rd_ptr_reg_46_ ( .D(n1847), .CLK(clk), .SN(1'b1), .Q(rd_ptr[46])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_47_ ( .D(n1787), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[47]) );
  DFFSNQ_X1 rd_ptr_reg_47_ ( .D(n1848), .CLK(clk), .SN(1'b1), .Q(rd_ptr[47])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_48_ ( .D(n1788), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[48]) );
  DFFSNQ_X1 rd_ptr_reg_48_ ( .D(n1849), .CLK(clk), .SN(1'b1), .Q(rd_ptr[48])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_49_ ( .D(n1789), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[49]) );
  DFFSNQ_X1 rd_ptr_reg_49_ ( .D(n1850), .CLK(clk), .SN(1'b1), .Q(rd_ptr[49])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_50_ ( .D(n1790), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[50]) );
  DFFSNQ_X1 rd_ptr_reg_50_ ( .D(n1851), .CLK(clk), .SN(1'b1), .Q(rd_ptr[50])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_51_ ( .D(n1791), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[51]) );
  DFFSNQ_X1 rd_ptr_reg_51_ ( .D(n1852), .CLK(clk), .SN(1'b1), .Q(rd_ptr[51])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_52_ ( .D(n1792), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[52]) );
  DFFSNQ_X1 rd_ptr_reg_52_ ( .D(n1853), .CLK(clk), .SN(1'b1), .Q(rd_ptr[52])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_53_ ( .D(n1793), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[53]) );
  DFFSNQ_X1 rd_ptr_reg_53_ ( .D(n1854), .CLK(clk), .SN(1'b1), .Q(rd_ptr[53])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_54_ ( .D(n1794), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[54]) );
  DFFSNQ_X1 rd_ptr_reg_54_ ( .D(n1855), .CLK(clk), .SN(1'b1), .Q(rd_ptr[54])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_55_ ( .D(n1795), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[55]) );
  DFFSNQ_X1 rd_ptr_reg_55_ ( .D(n1856), .CLK(clk), .SN(1'b1), .Q(rd_ptr[55])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_56_ ( .D(n1796), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[56]) );
  DFFSNQ_X1 rd_ptr_reg_56_ ( .D(n1857), .CLK(clk), .SN(1'b1), .Q(rd_ptr[56])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_57_ ( .D(n1797), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[57]) );
  DFFSNQ_X1 rd_ptr_reg_57_ ( .D(n1858), .CLK(clk), .SN(1'b1), .Q(rd_ptr[57])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_58_ ( .D(n1798), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[58]) );
  DFFSNQ_X1 rd_ptr_reg_58_ ( .D(n1859), .CLK(clk), .SN(1'b1), .Q(rd_ptr[58])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_59_ ( .D(n1799), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[59]) );
  DFFSNQ_X1 rd_ptr_reg_59_ ( .D(n1860), .CLK(clk), .SN(1'b1), .Q(rd_ptr[59])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_60_ ( .D(n1800), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[60]) );
  DFFSNQ_X1 rd_ptr_reg_60_ ( .D(n1861), .CLK(clk), .SN(1'b1), .Q(rd_ptr[60])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_61_ ( .D(n1801), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[61]) );
  DFFSNQ_X1 rd_ptr_reg_61_ ( .D(n1862), .CLK(clk), .SN(1'b1), .Q(rd_ptr[61])
         );
  DFFSNQ_X1 nxt_rd_ptr_reg_62_ ( .D(n1802), .CLK(clk), .SN(1'b1), .Q(
        nxt_rd_ptr[62]) );
  DFFSNQ_X1 rd_ptr_reg_62_ ( .D(n1863), .CLK(clk), .SN(1'b1), .Q(rd_ptr[62])
         );
  DFFSNQ_X1 rd_ptr_reg_63_ ( .D(n1864), .CLK(clk), .SN(1'b1), .Q(rd_ptr[63])
         );
  DFFSNQ_X1 full_reg ( .D(n1865), .CLK(clk), .SN(1'b1), .Q(full) );
  DFFSNQ_X1 wr_ptr_reg_0_ ( .D(n1866), .CLK(clk), .SN(1'b1), .Q(wr_ptr[0]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_1_ ( .D(n642), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[1]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_2_ ( .D(n641), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[2]) );
  DFFSNQ_X1 wr_ptr_reg_2_ ( .D(n948), .CLK(clk), .SN(1'b1), .Q(wr_ptr[2]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_3_ ( .D(n640), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[3]) );
  DFFSNQ_X1 wr_ptr_reg_3_ ( .D(n947), .CLK(clk), .SN(1'b1), .Q(wr_ptr[3]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_4_ ( .D(n639), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[4]) );
  DFFSNQ_X1 wr_ptr_reg_4_ ( .D(n1867), .CLK(clk), .SN(1'b1), .Q(wr_ptr[4]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_5_ ( .D(n638), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[5]) );
  DFFSNQ_X1 wr_ptr_reg_5_ ( .D(n946), .CLK(clk), .SN(1'b1), .Q(wr_ptr[5]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_6_ ( .D(n637), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[6]) );
  DFFSNQ_X1 wr_ptr_reg_6_ ( .D(n945), .CLK(clk), .SN(1'b1), .Q(wr_ptr[6]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_7_ ( .D(n636), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[7]) );
  DFFSNQ_X1 wr_ptr_reg_7_ ( .D(n944), .CLK(clk), .SN(1'b1), .Q(wr_ptr[7]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_8_ ( .D(n635), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[8]) );
  DFFSNQ_X1 wr_ptr_reg_8_ ( .D(n943), .CLK(clk), .SN(1'b1), .Q(wr_ptr[8]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_9_ ( .D(n634), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[9]) );
  DFFSNQ_X1 wr_ptr_reg_9_ ( .D(n942), .CLK(clk), .SN(1'b1), .Q(wr_ptr[9]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_10_ ( .D(n633), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[10]) );
  DFFSNQ_X1 wr_ptr_reg_10_ ( .D(n1868), .CLK(clk), .SN(1'b1), .Q(wr_ptr[10])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_11_ ( .D(n632), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[11]) );
  DFFSNQ_X1 wr_ptr_reg_11_ ( .D(n1869), .CLK(clk), .SN(1'b1), .Q(wr_ptr[11])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_12_ ( .D(n631), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[12]) );
  DFFSNQ_X1 wr_ptr_reg_12_ ( .D(n1870), .CLK(clk), .SN(1'b1), .Q(wr_ptr[12])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_13_ ( .D(n630), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[13]) );
  DFFSNQ_X1 wr_ptr_reg_13_ ( .D(n941), .CLK(clk), .SN(1'b1), .Q(wr_ptr[13]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_14_ ( .D(n629), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[14]) );
  DFFSNQ_X1 wr_ptr_reg_14_ ( .D(n940), .CLK(clk), .SN(1'b1), .Q(wr_ptr[14]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_15_ ( .D(n628), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[15]) );
  DFFSNQ_X1 wr_ptr_reg_15_ ( .D(n939), .CLK(clk), .SN(1'b1), .Q(wr_ptr[15]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_16_ ( .D(n627), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[16]) );
  DFFSNQ_X1 wr_ptr_reg_16_ ( .D(n938), .CLK(clk), .SN(1'b1), .Q(wr_ptr[16]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_17_ ( .D(n626), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[17]) );
  DFFSNQ_X1 wr_ptr_reg_17_ ( .D(n937), .CLK(clk), .SN(1'b1), .Q(wr_ptr[17]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_18_ ( .D(n625), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[18]) );
  DFFSNQ_X1 wr_ptr_reg_18_ ( .D(n936), .CLK(clk), .SN(1'b1), .Q(wr_ptr[18]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_19_ ( .D(n624), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[19]) );
  DFFSNQ_X1 wr_ptr_reg_19_ ( .D(n935), .CLK(clk), .SN(1'b1), .Q(wr_ptr[19]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_20_ ( .D(n623), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[20]) );
  DFFSNQ_X1 wr_ptr_reg_20_ ( .D(n934), .CLK(clk), .SN(1'b1), .Q(wr_ptr[20]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_21_ ( .D(n622), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[21]) );
  DFFSNQ_X1 wr_ptr_reg_21_ ( .D(n933), .CLK(clk), .SN(1'b1), .Q(wr_ptr[21]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_22_ ( .D(n621), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[22]) );
  DFFSNQ_X1 wr_ptr_reg_22_ ( .D(n932), .CLK(clk), .SN(1'b1), .Q(wr_ptr[22]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_23_ ( .D(n620), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[23]) );
  DFFSNQ_X1 wr_ptr_reg_23_ ( .D(n931), .CLK(clk), .SN(1'b1), .Q(wr_ptr[23]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_24_ ( .D(n619), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[24]) );
  DFFSNQ_X1 wr_ptr_reg_24_ ( .D(n930), .CLK(clk), .SN(1'b1), .Q(wr_ptr[24]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_25_ ( .D(n618), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[25]) );
  DFFSNQ_X1 wr_ptr_reg_25_ ( .D(n929), .CLK(clk), .SN(1'b1), .Q(wr_ptr[25]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_26_ ( .D(n617), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[26]) );
  DFFSNQ_X1 wr_ptr_reg_26_ ( .D(n928), .CLK(clk), .SN(1'b1), .Q(wr_ptr[26]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_27_ ( .D(n616), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[27]) );
  DFFSNQ_X1 wr_ptr_reg_27_ ( .D(n927), .CLK(clk), .SN(1'b1), .Q(wr_ptr[27]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_28_ ( .D(n615), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[28]) );
  DFFSNQ_X1 wr_ptr_reg_28_ ( .D(n926), .CLK(clk), .SN(1'b1), .Q(wr_ptr[28]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_29_ ( .D(n614), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[29]) );
  DFFSNQ_X1 wr_ptr_reg_29_ ( .D(n925), .CLK(clk), .SN(1'b1), .Q(wr_ptr[29]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_30_ ( .D(n613), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[30]) );
  DFFSNQ_X1 wr_ptr_reg_30_ ( .D(n924), .CLK(clk), .SN(1'b1), .Q(wr_ptr[30]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_31_ ( .D(n612), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[31]) );
  DFFSNQ_X1 wr_ptr_reg_31_ ( .D(n923), .CLK(clk), .SN(1'b1), .Q(wr_ptr[31]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_32_ ( .D(n611), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[32]) );
  DFFSNQ_X1 wr_ptr_reg_32_ ( .D(n922), .CLK(clk), .SN(1'b1), .Q(wr_ptr[32]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_33_ ( .D(n610), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[33]) );
  DFFSNQ_X1 wr_ptr_reg_33_ ( .D(n921), .CLK(clk), .SN(1'b1), .Q(wr_ptr[33]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_34_ ( .D(n609), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[34]) );
  DFFSNQ_X1 wr_ptr_reg_34_ ( .D(n920), .CLK(clk), .SN(1'b1), .Q(wr_ptr[34]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_35_ ( .D(n608), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[35]) );
  DFFSNQ_X1 wr_ptr_reg_35_ ( .D(n919), .CLK(clk), .SN(1'b1), .Q(wr_ptr[35]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_36_ ( .D(n607), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[36]) );
  DFFSNQ_X1 wr_ptr_reg_36_ ( .D(n918), .CLK(clk), .SN(1'b1), .Q(wr_ptr[36]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_37_ ( .D(n606), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[37]) );
  DFFSNQ_X1 wr_ptr_reg_37_ ( .D(n917), .CLK(clk), .SN(1'b1), .Q(wr_ptr[37]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_38_ ( .D(n605), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[38]) );
  DFFSNQ_X1 wr_ptr_reg_38_ ( .D(n916), .CLK(clk), .SN(1'b1), .Q(wr_ptr[38]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_39_ ( .D(n604), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[39]) );
  DFFSNQ_X1 wr_ptr_reg_39_ ( .D(n915), .CLK(clk), .SN(1'b1), .Q(wr_ptr[39]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_40_ ( .D(n603), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[40]) );
  DFFSNQ_X1 wr_ptr_reg_40_ ( .D(n914), .CLK(clk), .SN(1'b1), .Q(wr_ptr[40]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_41_ ( .D(n602), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[41]) );
  DFFSNQ_X1 wr_ptr_reg_41_ ( .D(n913), .CLK(clk), .SN(1'b1), .Q(wr_ptr[41]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_42_ ( .D(n601), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[42]) );
  DFFSNQ_X1 wr_ptr_reg_42_ ( .D(n912), .CLK(clk), .SN(1'b1), .Q(wr_ptr[42]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_43_ ( .D(n600), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[43]) );
  DFFSNQ_X1 wr_ptr_reg_43_ ( .D(n911), .CLK(clk), .SN(1'b1), .Q(wr_ptr[43]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_44_ ( .D(n599), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[44]) );
  DFFSNQ_X1 wr_ptr_reg_44_ ( .D(n910), .CLK(clk), .SN(1'b1), .Q(wr_ptr[44]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_45_ ( .D(n598), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[45]) );
  DFFSNQ_X1 wr_ptr_reg_45_ ( .D(n909), .CLK(clk), .SN(1'b1), .Q(wr_ptr[45]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_46_ ( .D(n597), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[46]) );
  DFFSNQ_X1 wr_ptr_reg_46_ ( .D(n1871), .CLK(clk), .SN(1'b1), .Q(wr_ptr[46])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_47_ ( .D(n596), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[47]) );
  DFFSNQ_X1 wr_ptr_reg_47_ ( .D(n1872), .CLK(clk), .SN(1'b1), .Q(wr_ptr[47])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_48_ ( .D(n595), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[48]) );
  DFFSNQ_X1 wr_ptr_reg_48_ ( .D(n1873), .CLK(clk), .SN(1'b1), .Q(wr_ptr[48])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_49_ ( .D(n594), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[49]) );
  DFFSNQ_X1 wr_ptr_reg_49_ ( .D(n1874), .CLK(clk), .SN(1'b1), .Q(wr_ptr[49])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_50_ ( .D(n593), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[50]) );
  DFFSNQ_X1 wr_ptr_reg_50_ ( .D(n1875), .CLK(clk), .SN(1'b1), .Q(wr_ptr[50])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_51_ ( .D(n592), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[51]) );
  DFFSNQ_X1 wr_ptr_reg_51_ ( .D(n1876), .CLK(clk), .SN(1'b1), .Q(wr_ptr[51])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_52_ ( .D(n591), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[52]) );
  DFFSNQ_X1 wr_ptr_reg_52_ ( .D(n1877), .CLK(clk), .SN(1'b1), .Q(wr_ptr[52])
         );
  DFFSNQ_X1 nxt_wr_ptr_reg_53_ ( .D(n590), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[53]) );
  DFFSNQ_X1 wr_ptr_reg_53_ ( .D(n908), .CLK(clk), .SN(1'b1), .Q(wr_ptr[53]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_54_ ( .D(n589), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[54]) );
  DFFSNQ_X1 wr_ptr_reg_54_ ( .D(n907), .CLK(clk), .SN(1'b1), .Q(wr_ptr[54]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_55_ ( .D(n588), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[55]) );
  DFFSNQ_X1 wr_ptr_reg_55_ ( .D(n906), .CLK(clk), .SN(1'b1), .Q(wr_ptr[55]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_56_ ( .D(n587), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[56]) );
  DFFSNQ_X1 wr_ptr_reg_56_ ( .D(n905), .CLK(clk), .SN(1'b1), .Q(wr_ptr[56]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_57_ ( .D(n586), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[57]) );
  DFFSNQ_X1 wr_ptr_reg_57_ ( .D(n904), .CLK(clk), .SN(1'b1), .Q(wr_ptr[57]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_58_ ( .D(n585), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[58]) );
  DFFSNQ_X1 wr_ptr_reg_58_ ( .D(n903), .CLK(clk), .SN(1'b1), .Q(wr_ptr[58]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_59_ ( .D(n584), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[59]) );
  DFFSNQ_X1 wr_ptr_reg_59_ ( .D(n902), .CLK(clk), .SN(1'b1), .Q(wr_ptr[59]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_60_ ( .D(n583), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[60]) );
  DFFSNQ_X1 wr_ptr_reg_60_ ( .D(n901), .CLK(clk), .SN(1'b1), .Q(wr_ptr[60]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_61_ ( .D(n582), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[61]) );
  DFFSNQ_X1 wr_ptr_reg_61_ ( .D(n900), .CLK(clk), .SN(1'b1), .Q(wr_ptr[61]) );
  DFFSNQ_X1 nxt_wr_ptr_reg_62_ ( .D(n581), .CLK(clk), .SN(1'b1), .Q(
        nxt_wr_ptr[62]) );
  DFFSNQ_X1 wr_ptr_reg_62_ ( .D(n899), .CLK(clk), .SN(1'b1), .Q(wr_ptr[62]) );
  DFFSNQ_X1 wr_ptr_reg_1_ ( .D(n949), .CLK(clk), .SN(1'b1), .Q(wr_ptr[1]) );
  DFFSNQ_X1 wr_ptr_reg_63_ ( .D(n644), .CLK(clk), .SN(1'b1), .Q(wr_ptr[63]) );
  DFFSNQ_X1 queue_reg_1__63_ ( .D(n1648), .CLK(clk), .SN(1'b1), .Q(queue[127])
         );
  DFFSNQ_X1 queue_reg_1__62_ ( .D(n1649), .CLK(clk), .SN(1'b1), .Q(queue[126])
         );
  DFFSNQ_X1 queue_reg_1__61_ ( .D(n1650), .CLK(clk), .SN(1'b1), .Q(queue[125])
         );
  DFFSNQ_X1 queue_reg_1__60_ ( .D(n1651), .CLK(clk), .SN(1'b1), .Q(queue[124])
         );
  DFFSNQ_X1 queue_reg_1__59_ ( .D(n1652), .CLK(clk), .SN(1'b1), .Q(queue[123])
         );
  DFFSNQ_X1 queue_reg_1__58_ ( .D(n1653), .CLK(clk), .SN(1'b1), .Q(queue[122])
         );
  DFFSNQ_X1 queue_reg_1__57_ ( .D(n1654), .CLK(clk), .SN(1'b1), .Q(queue[121])
         );
  DFFSNQ_X1 queue_reg_1__56_ ( .D(n1655), .CLK(clk), .SN(1'b1), .Q(queue[120])
         );
  DFFSNQ_X1 queue_reg_1__55_ ( .D(n1656), .CLK(clk), .SN(1'b1), .Q(queue[119])
         );
  DFFSNQ_X1 queue_reg_1__54_ ( .D(n1657), .CLK(clk), .SN(1'b1), .Q(queue[118])
         );
  DFFSNQ_X1 queue_reg_1__53_ ( .D(n1658), .CLK(clk), .SN(1'b1), .Q(queue[117])
         );
  DFFSNQ_X1 queue_reg_1__52_ ( .D(n1659), .CLK(clk), .SN(1'b1), .Q(queue[116])
         );
  DFFSNQ_X1 queue_reg_1__51_ ( .D(n1660), .CLK(clk), .SN(1'b1), .Q(queue[115])
         );
  DFFSNQ_X1 queue_reg_1__50_ ( .D(n1661), .CLK(clk), .SN(1'b1), .Q(queue[114])
         );
  DFFSNQ_X1 queue_reg_1__49_ ( .D(n1662), .CLK(clk), .SN(1'b1), .Q(queue[113])
         );
  DFFSNQ_X1 queue_reg_1__48_ ( .D(n1663), .CLK(clk), .SN(1'b1), .Q(queue[112])
         );
  DFFSNQ_X1 queue_reg_1__47_ ( .D(n1664), .CLK(clk), .SN(1'b1), .Q(queue[111])
         );
  DFFSNQ_X1 queue_reg_1__46_ ( .D(n1665), .CLK(clk), .SN(1'b1), .Q(queue[110])
         );
  DFFSNQ_X1 queue_reg_1__45_ ( .D(n1666), .CLK(clk), .SN(1'b1), .Q(queue[109])
         );
  DFFSNQ_X1 queue_reg_1__44_ ( .D(n1667), .CLK(clk), .SN(1'b1), .Q(queue[108])
         );
  DFFSNQ_X1 queue_reg_1__43_ ( .D(n1668), .CLK(clk), .SN(1'b1), .Q(queue[107])
         );
  DFFSNQ_X1 queue_reg_1__42_ ( .D(n1669), .CLK(clk), .SN(1'b1), .Q(queue[106])
         );
  DFFSNQ_X1 queue_reg_1__41_ ( .D(n1670), .CLK(clk), .SN(1'b1), .Q(queue[105])
         );
  DFFSNQ_X1 queue_reg_1__40_ ( .D(n1671), .CLK(clk), .SN(1'b1), .Q(queue[104])
         );
  DFFSNQ_X1 queue_reg_1__39_ ( .D(n1672), .CLK(clk), .SN(1'b1), .Q(queue[103])
         );
  DFFSNQ_X1 queue_reg_1__38_ ( .D(n1673), .CLK(clk), .SN(1'b1), .Q(queue[102])
         );
  DFFSNQ_X1 queue_reg_1__37_ ( .D(n1674), .CLK(clk), .SN(1'b1), .Q(queue[101])
         );
  DFFSNQ_X1 queue_reg_1__36_ ( .D(n1675), .CLK(clk), .SN(1'b1), .Q(queue[100])
         );
  DFFSNQ_X1 queue_reg_1__35_ ( .D(n1676), .CLK(clk), .SN(1'b1), .Q(queue[99])
         );
  DFFSNQ_X1 queue_reg_1__34_ ( .D(n1677), .CLK(clk), .SN(1'b1), .Q(queue[98])
         );
  DFFSNQ_X1 queue_reg_1__33_ ( .D(n1678), .CLK(clk), .SN(1'b1), .Q(queue[97])
         );
  DFFSNQ_X1 queue_reg_1__32_ ( .D(n1679), .CLK(clk), .SN(1'b1), .Q(queue[96])
         );
  DFFSNQ_X1 queue_reg_1__31_ ( .D(n1680), .CLK(clk), .SN(1'b1), .Q(queue[95])
         );
  DFFSNQ_X1 queue_reg_1__30_ ( .D(n1681), .CLK(clk), .SN(1'b1), .Q(queue[94])
         );
  DFFSNQ_X1 queue_reg_1__29_ ( .D(n1682), .CLK(clk), .SN(1'b1), .Q(queue[93])
         );
  DFFSNQ_X1 queue_reg_1__28_ ( .D(n1683), .CLK(clk), .SN(1'b1), .Q(queue[92])
         );
  DFFSNQ_X1 queue_reg_1__27_ ( .D(n1684), .CLK(clk), .SN(1'b1), .Q(queue[91])
         );
  DFFSNQ_X1 queue_reg_1__26_ ( .D(n1685), .CLK(clk), .SN(1'b1), .Q(queue[90])
         );
  DFFSNQ_X1 queue_reg_1__25_ ( .D(n1686), .CLK(clk), .SN(1'b1), .Q(queue[89])
         );
  DFFSNQ_X1 queue_reg_1__24_ ( .D(n1687), .CLK(clk), .SN(1'b1), .Q(queue[88])
         );
  DFFSNQ_X1 queue_reg_1__23_ ( .D(n1688), .CLK(clk), .SN(1'b1), .Q(queue[87])
         );
  DFFSNQ_X1 queue_reg_1__22_ ( .D(n1689), .CLK(clk), .SN(1'b1), .Q(queue[86])
         );
  DFFSNQ_X1 queue_reg_1__21_ ( .D(n1690), .CLK(clk), .SN(1'b1), .Q(queue[85])
         );
  DFFSNQ_X1 queue_reg_1__20_ ( .D(n1691), .CLK(clk), .SN(1'b1), .Q(queue[84])
         );
  DFFSNQ_X1 queue_reg_1__19_ ( .D(n1692), .CLK(clk), .SN(1'b1), .Q(queue[83])
         );
  DFFSNQ_X1 queue_reg_1__18_ ( .D(n1693), .CLK(clk), .SN(1'b1), .Q(queue[82])
         );
  DFFSNQ_X1 queue_reg_1__17_ ( .D(n1694), .CLK(clk), .SN(1'b1), .Q(queue[81])
         );
  DFFSNQ_X1 queue_reg_1__16_ ( .D(n1695), .CLK(clk), .SN(1'b1), .Q(queue[80])
         );
  DFFSNQ_X1 queue_reg_1__15_ ( .D(n1696), .CLK(clk), .SN(1'b1), .Q(queue[79])
         );
  DFFSNQ_X1 queue_reg_1__14_ ( .D(n1697), .CLK(clk), .SN(1'b1), .Q(queue[78])
         );
  DFFSNQ_X1 queue_reg_1__13_ ( .D(n1698), .CLK(clk), .SN(1'b1), .Q(queue[77])
         );
  DFFSNQ_X1 queue_reg_1__12_ ( .D(n1699), .CLK(clk), .SN(1'b1), .Q(queue[76])
         );
  DFFSNQ_X1 queue_reg_1__11_ ( .D(n1700), .CLK(clk), .SN(1'b1), .Q(queue[75])
         );
  DFFSNQ_X1 queue_reg_1__10_ ( .D(n1701), .CLK(clk), .SN(1'b1), .Q(queue[74])
         );
  DFFSNQ_X1 queue_reg_1__9_ ( .D(n1702), .CLK(clk), .SN(1'b1), .Q(queue[73])
         );
  DFFSNQ_X1 queue_reg_1__8_ ( .D(n1703), .CLK(clk), .SN(1'b1), .Q(queue[72])
         );
  DFFSNQ_X1 queue_reg_1__7_ ( .D(n1704), .CLK(clk), .SN(1'b1), .Q(queue[71])
         );
  DFFSNQ_X1 queue_reg_1__6_ ( .D(n1705), .CLK(clk), .SN(1'b1), .Q(queue[70])
         );
  DFFSNQ_X1 queue_reg_1__5_ ( .D(n1706), .CLK(clk), .SN(1'b1), .Q(queue[69])
         );
  DFFSNQ_X1 queue_reg_1__4_ ( .D(n1707), .CLK(clk), .SN(1'b1), .Q(queue[68])
         );
  DFFSNQ_X1 queue_reg_1__3_ ( .D(n1708), .CLK(clk), .SN(1'b1), .Q(queue[67])
         );
  DFFSNQ_X1 queue_reg_1__2_ ( .D(n1709), .CLK(clk), .SN(1'b1), .Q(queue[66])
         );
  DFFSNQ_X1 queue_reg_1__1_ ( .D(n1710), .CLK(clk), .SN(1'b1), .Q(queue[65])
         );
  DFFSNQ_X1 queue_reg_1__0_ ( .D(n1711), .CLK(clk), .SN(1'b1), .Q(queue[64])
         );
  DFFSNQ_X1 queue_reg_0__63_ ( .D(n951), .CLK(clk), .SN(1'b1), .Q(queue[63])
         );
  DFFSNQ_X1 queue_reg_0__62_ ( .D(n952), .CLK(clk), .SN(1'b1), .Q(queue[62])
         );
  DFFSNQ_X1 queue_reg_0__61_ ( .D(n953), .CLK(clk), .SN(1'b1), .Q(queue[61])
         );
  DFFSNQ_X1 queue_reg_0__60_ ( .D(n954), .CLK(clk), .SN(1'b1), .Q(queue[60])
         );
  DFFSNQ_X1 queue_reg_0__59_ ( .D(n955), .CLK(clk), .SN(1'b1), .Q(queue[59])
         );
  DFFSNQ_X1 queue_reg_0__58_ ( .D(n956), .CLK(clk), .SN(1'b1), .Q(queue[58])
         );
  DFFSNQ_X1 queue_reg_0__57_ ( .D(n957), .CLK(clk), .SN(1'b1), .Q(queue[57])
         );
  DFFSNQ_X1 queue_reg_0__56_ ( .D(n958), .CLK(clk), .SN(1'b1), .Q(queue[56])
         );
  DFFSNQ_X1 queue_reg_0__55_ ( .D(n959), .CLK(clk), .SN(1'b1), .Q(queue[55])
         );
  DFFSNQ_X1 queue_reg_0__54_ ( .D(n960), .CLK(clk), .SN(1'b1), .Q(queue[54])
         );
  DFFSNQ_X1 queue_reg_0__53_ ( .D(n961), .CLK(clk), .SN(1'b1), .Q(queue[53])
         );
  DFFSNQ_X1 queue_reg_0__52_ ( .D(n962), .CLK(clk), .SN(1'b1), .Q(queue[52])
         );
  DFFSNQ_X1 queue_reg_0__51_ ( .D(n963), .CLK(clk), .SN(1'b1), .Q(queue[51])
         );
  DFFSNQ_X1 queue_reg_0__50_ ( .D(n964), .CLK(clk), .SN(1'b1), .Q(queue[50])
         );
  DFFSNQ_X1 queue_reg_0__49_ ( .D(n965), .CLK(clk), .SN(1'b1), .Q(queue[49])
         );
  DFFSNQ_X1 queue_reg_0__48_ ( .D(n966), .CLK(clk), .SN(1'b1), .Q(queue[48])
         );
  DFFSNQ_X1 queue_reg_0__47_ ( .D(n967), .CLK(clk), .SN(1'b1), .Q(queue[47])
         );
  DFFSNQ_X1 queue_reg_0__46_ ( .D(n968), .CLK(clk), .SN(1'b1), .Q(queue[46])
         );
  DFFSNQ_X1 queue_reg_0__45_ ( .D(n969), .CLK(clk), .SN(1'b1), .Q(queue[45])
         );
  DFFSNQ_X1 queue_reg_0__44_ ( .D(n970), .CLK(clk), .SN(1'b1), .Q(queue[44])
         );
  DFFSNQ_X1 queue_reg_0__43_ ( .D(n971), .CLK(clk), .SN(1'b1), .Q(queue[43])
         );
  DFFSNQ_X1 queue_reg_0__42_ ( .D(n972), .CLK(clk), .SN(1'b1), .Q(queue[42])
         );
  DFFSNQ_X1 queue_reg_0__41_ ( .D(n973), .CLK(clk), .SN(1'b1), .Q(queue[41])
         );
  DFFSNQ_X1 queue_reg_0__40_ ( .D(n974), .CLK(clk), .SN(1'b1), .Q(queue[40])
         );
  DFFSNQ_X1 queue_reg_0__39_ ( .D(n975), .CLK(clk), .SN(1'b1), .Q(queue[39])
         );
  DFFSNQ_X1 queue_reg_0__38_ ( .D(n976), .CLK(clk), .SN(1'b1), .Q(queue[38])
         );
  DFFSNQ_X1 queue_reg_0__37_ ( .D(n1336), .CLK(clk), .SN(1'b1), .Q(queue[37])
         );
  DFFSNQ_X1 queue_reg_0__36_ ( .D(n1611), .CLK(clk), .SN(1'b1), .Q(queue[36])
         );
  DFFSNQ_X1 queue_reg_0__35_ ( .D(n1612), .CLK(clk), .SN(1'b1), .Q(queue[35])
         );
  DFFSNQ_X1 queue_reg_0__34_ ( .D(n1613), .CLK(clk), .SN(1'b1), .Q(queue[34])
         );
  DFFSNQ_X1 queue_reg_0__33_ ( .D(n1614), .CLK(clk), .SN(1'b1), .Q(queue[33])
         );
  DFFSNQ_X1 queue_reg_0__32_ ( .D(n1615), .CLK(clk), .SN(1'b1), .Q(queue[32])
         );
  DFFSNQ_X1 queue_reg_0__31_ ( .D(n1616), .CLK(clk), .SN(1'b1), .Q(queue[31])
         );
  DFFSNQ_X1 queue_reg_0__30_ ( .D(n1617), .CLK(clk), .SN(1'b1), .Q(queue[30])
         );
  DFFSNQ_X1 queue_reg_0__29_ ( .D(n1618), .CLK(clk), .SN(1'b1), .Q(queue[29])
         );
  DFFSNQ_X1 queue_reg_0__28_ ( .D(n1619), .CLK(clk), .SN(1'b1), .Q(queue[28])
         );
  DFFSNQ_X1 queue_reg_0__27_ ( .D(n1620), .CLK(clk), .SN(1'b1), .Q(queue[27])
         );
  DFFSNQ_X1 queue_reg_0__26_ ( .D(n1621), .CLK(clk), .SN(1'b1), .Q(queue[26])
         );
  DFFSNQ_X1 queue_reg_0__25_ ( .D(n1622), .CLK(clk), .SN(1'b1), .Q(queue[25])
         );
  DFFSNQ_X1 queue_reg_0__24_ ( .D(n1623), .CLK(clk), .SN(1'b1), .Q(queue[24])
         );
  DFFSNQ_X1 queue_reg_0__23_ ( .D(n1624), .CLK(clk), .SN(1'b1), .Q(queue[23])
         );
  DFFSNQ_X1 queue_reg_0__22_ ( .D(n1625), .CLK(clk), .SN(1'b1), .Q(queue[22])
         );
  DFFSNQ_X1 queue_reg_0__21_ ( .D(n1626), .CLK(clk), .SN(1'b1), .Q(queue[21])
         );
  DFFSNQ_X1 queue_reg_0__20_ ( .D(n1627), .CLK(clk), .SN(1'b1), .Q(queue[20])
         );
  DFFSNQ_X1 queue_reg_0__19_ ( .D(n1628), .CLK(clk), .SN(1'b1), .Q(queue[19])
         );
  DFFSNQ_X1 queue_reg_0__18_ ( .D(n1629), .CLK(clk), .SN(1'b1), .Q(queue[18])
         );
  DFFSNQ_X1 queue_reg_0__17_ ( .D(n1630), .CLK(clk), .SN(1'b1), .Q(queue[17])
         );
  DFFSNQ_X1 queue_reg_0__16_ ( .D(n1631), .CLK(clk), .SN(1'b1), .Q(queue[16])
         );
  DFFSNQ_X1 queue_reg_0__15_ ( .D(n1632), .CLK(clk), .SN(1'b1), .Q(queue[15])
         );
  DFFSNQ_X1 queue_reg_0__14_ ( .D(n1633), .CLK(clk), .SN(1'b1), .Q(queue[14])
         );
  DFFSNQ_X1 queue_reg_0__13_ ( .D(n1634), .CLK(clk), .SN(1'b1), .Q(queue[13])
         );
  DFFSNQ_X1 queue_reg_0__12_ ( .D(n1635), .CLK(clk), .SN(1'b1), .Q(queue[12])
         );
  DFFSNQ_X1 queue_reg_0__11_ ( .D(n1636), .CLK(clk), .SN(1'b1), .Q(queue[11])
         );
  DFFSNQ_X1 queue_reg_0__10_ ( .D(n1637), .CLK(clk), .SN(1'b1), .Q(queue[10])
         );
  DFFSNQ_X1 queue_reg_0__9_ ( .D(n1638), .CLK(clk), .SN(1'b1), .Q(queue[9]) );
  DFFSNQ_X1 queue_reg_0__8_ ( .D(n1639), .CLK(clk), .SN(1'b1), .Q(queue[8]) );
  DFFSNQ_X1 queue_reg_0__7_ ( .D(n1640), .CLK(clk), .SN(1'b1), .Q(queue[7]) );
  DFFSNQ_X1 queue_reg_0__6_ ( .D(n1641), .CLK(clk), .SN(1'b1), .Q(queue[6]) );
  DFFSNQ_X1 queue_reg_0__5_ ( .D(n1642), .CLK(clk), .SN(1'b1), .Q(queue[5]) );
  DFFSNQ_X1 queue_reg_0__4_ ( .D(n1643), .CLK(clk), .SN(1'b1), .Q(queue[4]) );
  DFFSNQ_X1 queue_reg_0__3_ ( .D(n1644), .CLK(clk), .SN(1'b1), .Q(queue[3]) );
  DFFSNQ_X1 queue_reg_0__2_ ( .D(n1645), .CLK(clk), .SN(1'b1), .Q(queue[2]) );
  DFFSNQ_X1 queue_reg_0__1_ ( .D(n1646), .CLK(clk), .SN(1'b1), .Q(queue[1]) );
  DFFSNQ_X1 queue_reg_0__0_ ( .D(n1647), .CLK(clk), .SN(1'b1), .Q(queue[0]) );
  DFFSNQ_X1 data_out_reg_63_ ( .D(n645), .CLK(clk), .SN(1'b1), .Q(data_out[63]) );
  DFFSNQ_X1 data_out_reg_62_ ( .D(n646), .CLK(clk), .SN(1'b1), .Q(data_out[62]) );
  DFFSNQ_X1 data_out_reg_61_ ( .D(n647), .CLK(clk), .SN(1'b1), .Q(data_out[61]) );
  DFFSNQ_X1 data_out_reg_60_ ( .D(n648), .CLK(clk), .SN(1'b1), .Q(data_out[60]) );
  DFFSNQ_X1 data_out_reg_59_ ( .D(n649), .CLK(clk), .SN(1'b1), .Q(data_out[59]) );
  DFFSNQ_X1 data_out_reg_58_ ( .D(n650), .CLK(clk), .SN(1'b1), .Q(data_out[58]) );
  DFFSNQ_X1 data_out_reg_57_ ( .D(n651), .CLK(clk), .SN(1'b1), .Q(data_out[57]) );
  DFFSNQ_X1 data_out_reg_56_ ( .D(n652), .CLK(clk), .SN(1'b1), .Q(data_out[56]) );
  DFFSNQ_X1 data_out_reg_55_ ( .D(n653), .CLK(clk), .SN(1'b1), .Q(data_out[55]) );
  DFFSNQ_X1 data_out_reg_54_ ( .D(n654), .CLK(clk), .SN(1'b1), .Q(data_out[54]) );
  DFFSNQ_X1 data_out_reg_53_ ( .D(n655), .CLK(clk), .SN(1'b1), .Q(data_out[53]) );
  DFFSNQ_X1 data_out_reg_52_ ( .D(n656), .CLK(clk), .SN(1'b1), .Q(data_out[52]) );
  DFFSNQ_X1 data_out_reg_51_ ( .D(n657), .CLK(clk), .SN(1'b1), .Q(data_out[51]) );
  DFFSNQ_X1 data_out_reg_50_ ( .D(n658), .CLK(clk), .SN(1'b1), .Q(data_out[50]) );
  DFFSNQ_X1 data_out_reg_49_ ( .D(n659), .CLK(clk), .SN(1'b1), .Q(data_out[49]) );
  DFFSNQ_X1 data_out_reg_48_ ( .D(n660), .CLK(clk), .SN(1'b1), .Q(data_out[48]) );
  DFFSNQ_X1 data_out_reg_47_ ( .D(n661), .CLK(clk), .SN(1'b1), .Q(data_out[47]) );
  DFFSNQ_X1 data_out_reg_46_ ( .D(n662), .CLK(clk), .SN(1'b1), .Q(data_out[46]) );
  DFFSNQ_X1 data_out_reg_45_ ( .D(n663), .CLK(clk), .SN(1'b1), .Q(data_out[45]) );
  DFFSNQ_X1 data_out_reg_44_ ( .D(n664), .CLK(clk), .SN(1'b1), .Q(data_out[44]) );
  DFFSNQ_X1 data_out_reg_43_ ( .D(n665), .CLK(clk), .SN(1'b1), .Q(data_out[43]) );
  DFFSNQ_X1 data_out_reg_42_ ( .D(n666), .CLK(clk), .SN(1'b1), .Q(data_out[42]) );
  DFFSNQ_X1 data_out_reg_41_ ( .D(n667), .CLK(clk), .SN(1'b1), .Q(data_out[41]) );
  DFFSNQ_X1 data_out_reg_40_ ( .D(n668), .CLK(clk), .SN(1'b1), .Q(data_out[40]) );
  DFFSNQ_X1 data_out_reg_39_ ( .D(n669), .CLK(clk), .SN(1'b1), .Q(data_out[39]) );
  DFFSNQ_X1 data_out_reg_38_ ( .D(n670), .CLK(clk), .SN(1'b1), .Q(data_out[38]) );
  DFFSNQ_X1 data_out_reg_37_ ( .D(n671), .CLK(clk), .SN(1'b1), .Q(data_out[37]) );
  DFFSNQ_X1 data_out_reg_36_ ( .D(n672), .CLK(clk), .SN(1'b1), .Q(data_out[36]) );
  DFFSNQ_X1 data_out_reg_35_ ( .D(n673), .CLK(clk), .SN(1'b1), .Q(data_out[35]) );
  DFFSNQ_X1 data_out_reg_34_ ( .D(n674), .CLK(clk), .SN(1'b1), .Q(data_out[34]) );
  DFFSNQ_X1 data_out_reg_33_ ( .D(n675), .CLK(clk), .SN(1'b1), .Q(data_out[33]) );
  DFFSNQ_X1 data_out_reg_32_ ( .D(n676), .CLK(clk), .SN(1'b1), .Q(data_out[32]) );
  DFFSNQ_X1 data_out_reg_31_ ( .D(n677), .CLK(clk), .SN(1'b1), .Q(data_out[31]) );
  DFFSNQ_X1 data_out_reg_30_ ( .D(n678), .CLK(clk), .SN(1'b1), .Q(data_out[30]) );
  DFFSNQ_X1 data_out_reg_29_ ( .D(n679), .CLK(clk), .SN(1'b1), .Q(data_out[29]) );
  DFFSNQ_X1 data_out_reg_28_ ( .D(n680), .CLK(clk), .SN(1'b1), .Q(data_out[28]) );
  DFFSNQ_X1 data_out_reg_27_ ( .D(n681), .CLK(clk), .SN(1'b1), .Q(data_out[27]) );
  DFFSNQ_X1 data_out_reg_26_ ( .D(n682), .CLK(clk), .SN(1'b1), .Q(data_out[26]) );
  DFFSNQ_X1 data_out_reg_25_ ( .D(n683), .CLK(clk), .SN(1'b1), .Q(data_out[25]) );
  DFFSNQ_X1 data_out_reg_24_ ( .D(n684), .CLK(clk), .SN(1'b1), .Q(data_out[24]) );
  DFFSNQ_X1 data_out_reg_23_ ( .D(n685), .CLK(clk), .SN(1'b1), .Q(data_out[23]) );
  DFFSNQ_X1 data_out_reg_22_ ( .D(n686), .CLK(clk), .SN(1'b1), .Q(data_out[22]) );
  DFFSNQ_X1 data_out_reg_21_ ( .D(n687), .CLK(clk), .SN(1'b1), .Q(data_out[21]) );
  DFFSNQ_X1 data_out_reg_20_ ( .D(n688), .CLK(clk), .SN(1'b1), .Q(data_out[20]) );
  DFFSNQ_X1 data_out_reg_19_ ( .D(n689), .CLK(clk), .SN(1'b1), .Q(data_out[19]) );
  DFFSNQ_X1 data_out_reg_18_ ( .D(n690), .CLK(clk), .SN(1'b1), .Q(data_out[18]) );
  DFFSNQ_X1 data_out_reg_17_ ( .D(n691), .CLK(clk), .SN(1'b1), .Q(data_out[17]) );
  DFFSNQ_X1 data_out_reg_16_ ( .D(n692), .CLK(clk), .SN(1'b1), .Q(data_out[16]) );
  DFFSNQ_X1 data_out_reg_15_ ( .D(n693), .CLK(clk), .SN(1'b1), .Q(data_out[15]) );
  DFFSNQ_X1 data_out_reg_14_ ( .D(n694), .CLK(clk), .SN(1'b1), .Q(data_out[14]) );
  DFFSNQ_X1 data_out_reg_13_ ( .D(n695), .CLK(clk), .SN(1'b1), .Q(data_out[13]) );
  DFFSNQ_X1 data_out_reg_12_ ( .D(n696), .CLK(clk), .SN(1'b1), .Q(data_out[12]) );
  DFFSNQ_X1 data_out_reg_11_ ( .D(n697), .CLK(clk), .SN(1'b1), .Q(data_out[11]) );
  DFFSNQ_X1 data_out_reg_10_ ( .D(n698), .CLK(clk), .SN(1'b1), .Q(data_out[10]) );
  DFFSNQ_X1 data_out_reg_9_ ( .D(n699), .CLK(clk), .SN(1'b1), .Q(data_out[9])
         );
  DFFSNQ_X1 data_out_reg_8_ ( .D(n700), .CLK(clk), .SN(1'b1), .Q(data_out[8])
         );
  DFFSNQ_X1 data_out_reg_7_ ( .D(n701), .CLK(clk), .SN(1'b1), .Q(data_out[7])
         );
  DFFSNQ_X1 data_out_reg_6_ ( .D(n702), .CLK(clk), .SN(1'b1), .Q(data_out[6])
         );
  DFFSNQ_X1 data_out_reg_5_ ( .D(n703), .CLK(clk), .SN(1'b1), .Q(data_out[5])
         );
  DFFSNQ_X1 data_out_reg_4_ ( .D(n704), .CLK(clk), .SN(1'b1), .Q(data_out[4])
         );
  DFFSNQ_X1 data_out_reg_3_ ( .D(n705), .CLK(clk), .SN(1'b1), .Q(data_out[3])
         );
  DFFSNQ_X1 data_out_reg_2_ ( .D(n706), .CLK(clk), .SN(1'b1), .Q(data_out[2])
         );
  DFFSNQ_X1 data_out_reg_1_ ( .D(n707), .CLK(clk), .SN(1'b1), .Q(data_out[1])
         );
  DFFSNQ_X1 data_out_reg_0_ ( .D(n708), .CLK(clk), .SN(1'b1), .Q(data_out[0])
         );
  AND2_X1 U1528 ( .A1(n1736), .A2(n2303), .Z(n2367) );
  AND2_X1 U1529 ( .A1(n2148), .A2(n2147), .Z(n2217) );
  OR4_X1 U1530 ( .A1(wr_ptr[40]), .A2(wr_ptr[41]), .A3(wr_ptr[3]), .A4(n2142), 
        .Z(n2145) );
  OR4_X1 U1531 ( .A1(wr_ptr[45]), .A2(wr_ptr[44]), .A3(wr_ptr[43]), .A4(
        wr_ptr[42]), .Z(n2142) );
  OR4_X1 U1532 ( .A1(wr_ptr[17]), .A2(wr_ptr[18]), .A3(wr_ptr[19]), .A4(
        wr_ptr[20]), .Z(n2134) );
  OR4_X1 U1533 ( .A1(wr_ptr[21]), .A2(wr_ptr[22]), .A3(wr_ptr[23]), .A4(
        wr_ptr[24]), .Z(n2135) );
  AND2_X1 U1534 ( .A1(n2011), .A2(n1736), .Z(n1985) );
  XOR2_X1 U1535 ( .A1(n874), .A2(nxt_wr_ptr[51]), .Z(n1973) );
  XOR2_X1 U1536 ( .A1(n872), .A2(nxt_wr_ptr[50]), .Z(n1974) );
  XOR2_X1 U1537 ( .A1(n870), .A2(nxt_wr_ptr[49]), .Z(n1975) );
  XOR2_X1 U1538 ( .A1(n868), .A2(nxt_wr_ptr[48]), .Z(n1976) );
  XOR2_X1 U1539 ( .A1(n882), .A2(nxt_wr_ptr[55]), .Z(n1969) );
  XOR2_X1 U1540 ( .A1(n880), .A2(nxt_wr_ptr[54]), .Z(n1970) );
  XOR2_X1 U1541 ( .A1(n878), .A2(nxt_wr_ptr[53]), .Z(n1971) );
  XOR2_X1 U1542 ( .A1(n876), .A2(nxt_wr_ptr[52]), .Z(n1972) );
  XOR2_X1 U1543 ( .A1(n890), .A2(nxt_wr_ptr[59]), .Z(n1965) );
  XOR2_X1 U1544 ( .A1(n888), .A2(nxt_wr_ptr[58]), .Z(n1966) );
  XOR2_X1 U1545 ( .A1(n886), .A2(nxt_wr_ptr[57]), .Z(n1967) );
  XOR2_X1 U1546 ( .A1(n884), .A2(nxt_wr_ptr[56]), .Z(n1968) );
  XOR2_X1 U1547 ( .A1(n775), .A2(nxt_wr_ptr[63]), .Z(n1961) );
  XOR2_X1 U1548 ( .A1(n896), .A2(nxt_wr_ptr[62]), .Z(n1962) );
  XOR2_X1 U1549 ( .A1(n894), .A2(nxt_wr_ptr[61]), .Z(n1963) );
  XOR2_X1 U1550 ( .A1(n892), .A2(nxt_wr_ptr[60]), .Z(n1964) );
  XOR2_X1 U1551 ( .A1(n842), .A2(nxt_wr_ptr[35]), .Z(n1953) );
  XOR2_X1 U1552 ( .A1(n840), .A2(nxt_wr_ptr[34]), .Z(n1954) );
  XOR2_X1 U1553 ( .A1(n838), .A2(nxt_wr_ptr[33]), .Z(n1955) );
  XOR2_X1 U1554 ( .A1(n836), .A2(nxt_wr_ptr[32]), .Z(n1956) );
  XOR2_X1 U1555 ( .A1(n850), .A2(nxt_wr_ptr[39]), .Z(n1949) );
  XOR2_X1 U1556 ( .A1(n848), .A2(nxt_wr_ptr[38]), .Z(n1950) );
  XOR2_X1 U1557 ( .A1(n846), .A2(nxt_wr_ptr[37]), .Z(n1951) );
  XOR2_X1 U1558 ( .A1(n844), .A2(nxt_wr_ptr[36]), .Z(n1952) );
  XOR2_X1 U1559 ( .A1(n858), .A2(nxt_wr_ptr[43]), .Z(n1945) );
  XOR2_X1 U1560 ( .A1(n856), .A2(nxt_wr_ptr[42]), .Z(n1946) );
  XOR2_X1 U1561 ( .A1(n854), .A2(nxt_wr_ptr[41]), .Z(n1947) );
  XOR2_X1 U1562 ( .A1(n852), .A2(nxt_wr_ptr[40]), .Z(n1948) );
  XOR2_X1 U1563 ( .A1(n866), .A2(nxt_wr_ptr[47]), .Z(n1941) );
  XOR2_X1 U1564 ( .A1(n864), .A2(nxt_wr_ptr[46]), .Z(n1942) );
  XOR2_X1 U1565 ( .A1(n862), .A2(nxt_wr_ptr[45]), .Z(n1943) );
  XOR2_X1 U1566 ( .A1(n860), .A2(nxt_wr_ptr[44]), .Z(n1944) );
  XOR2_X1 U1567 ( .A1(n810), .A2(nxt_wr_ptr[19]), .Z(n1933) );
  XOR2_X1 U1568 ( .A1(n808), .A2(nxt_wr_ptr[18]), .Z(n1934) );
  XOR2_X1 U1569 ( .A1(n806), .A2(nxt_wr_ptr[17]), .Z(n1935) );
  XOR2_X1 U1570 ( .A1(n804), .A2(nxt_wr_ptr[16]), .Z(n1936) );
  XOR2_X1 U1571 ( .A1(n818), .A2(nxt_wr_ptr[23]), .Z(n1929) );
  XOR2_X1 U1572 ( .A1(n816), .A2(nxt_wr_ptr[22]), .Z(n1930) );
  XOR2_X1 U1573 ( .A1(n814), .A2(nxt_wr_ptr[21]), .Z(n1931) );
  XOR2_X1 U1574 ( .A1(n812), .A2(nxt_wr_ptr[20]), .Z(n1932) );
  XOR2_X1 U1575 ( .A1(n826), .A2(nxt_wr_ptr[27]), .Z(n1925) );
  XOR2_X1 U1576 ( .A1(n824), .A2(nxt_wr_ptr[26]), .Z(n1926) );
  XOR2_X1 U1577 ( .A1(n822), .A2(nxt_wr_ptr[25]), .Z(n1927) );
  XOR2_X1 U1578 ( .A1(n820), .A2(nxt_wr_ptr[24]), .Z(n1928) );
  XOR2_X1 U1579 ( .A1(n834), .A2(nxt_wr_ptr[31]), .Z(n1921) );
  XOR2_X1 U1580 ( .A1(n832), .A2(nxt_wr_ptr[30]), .Z(n1922) );
  XOR2_X1 U1581 ( .A1(n830), .A2(nxt_wr_ptr[29]), .Z(n1923) );
  XOR2_X1 U1582 ( .A1(n828), .A2(nxt_wr_ptr[28]), .Z(n1924) );
  XOR2_X1 U1583 ( .A1(n778), .A2(nxt_wr_ptr[3]), .Z(n1913) );
  XOR2_X1 U1584 ( .A1(n777), .A2(nxt_wr_ptr[2]), .Z(n1914) );
  XOR2_X1 U1585 ( .A1(n776), .A2(nxt_wr_ptr[1]), .Z(n1915) );
  XOR2_X1 U1586 ( .A1(n774), .A2(nxt_wr_ptr[0]), .Z(n1916) );
  XOR2_X1 U1587 ( .A1(n786), .A2(nxt_wr_ptr[7]), .Z(n1909) );
  XOR2_X1 U1588 ( .A1(n784), .A2(nxt_wr_ptr[6]), .Z(n1910) );
  XOR2_X1 U1589 ( .A1(n782), .A2(nxt_wr_ptr[5]), .Z(n1911) );
  XOR2_X1 U1590 ( .A1(n780), .A2(nxt_wr_ptr[4]), .Z(n1912) );
  XOR2_X1 U1591 ( .A1(n794), .A2(nxt_wr_ptr[11]), .Z(n1905) );
  XOR2_X1 U1592 ( .A1(n792), .A2(nxt_wr_ptr[10]), .Z(n1906) );
  XOR2_X1 U1593 ( .A1(n790), .A2(nxt_wr_ptr[9]), .Z(n1907) );
  XOR2_X1 U1594 ( .A1(n788), .A2(nxt_wr_ptr[8]), .Z(n1908) );
  XOR2_X1 U1595 ( .A1(n802), .A2(nxt_wr_ptr[15]), .Z(n1901) );
  XOR2_X1 U1596 ( .A1(n800), .A2(nxt_wr_ptr[14]), .Z(n1902) );
  XOR2_X1 U1597 ( .A1(n798), .A2(nxt_wr_ptr[13]), .Z(n1903) );
  XOR2_X1 U1598 ( .A1(n796), .A2(nxt_wr_ptr[12]), .Z(n1904) );
  AND2_X1 U1599 ( .A1(n471), .A2(n1899), .Z(n2073) );
  OR4_X1 U1600 ( .A1(nxt_wr_ptr[53]), .A2(nxt_wr_ptr[54]), .A3(nxt_wr_ptr[55]), 
        .A4(nxt_wr_ptr[56]), .Z(n1890) );
  OR4_X1 U1601 ( .A1(nxt_wr_ptr[57]), .A2(nxt_wr_ptr[58]), .A3(nxt_wr_ptr[59]), 
        .A4(nxt_wr_ptr[5]), .Z(n1891) );
  OR4_X1 U1602 ( .A1(nxt_wr_ptr[60]), .A2(nxt_wr_ptr[61]), .A3(nxt_wr_ptr[62]), 
        .A4(nxt_wr_ptr[63]), .Z(n1892) );
  OR4_X1 U1603 ( .A1(nxt_wr_ptr[6]), .A2(nxt_wr_ptr[7]), .A3(nxt_wr_ptr[8]), 
        .A4(nxt_wr_ptr[9]), .Z(n1893) );
  OR4_X1 U1604 ( .A1(nxt_wr_ptr[39]), .A2(nxt_wr_ptr[3]), .A3(nxt_wr_ptr[40]), 
        .A4(nxt_wr_ptr[41]), .Z(n1886) );
  OR4_X1 U1605 ( .A1(nxt_wr_ptr[42]), .A2(nxt_wr_ptr[43]), .A3(nxt_wr_ptr[44]), 
        .A4(nxt_wr_ptr[45]), .Z(n1887) );
  OR4_X1 U1606 ( .A1(nxt_wr_ptr[24]), .A2(nxt_wr_ptr[25]), .A3(nxt_wr_ptr[26]), 
        .A4(nxt_wr_ptr[27]), .Z(n1882) );
  OR4_X1 U1607 ( .A1(nxt_wr_ptr[28]), .A2(nxt_wr_ptr[29]), .A3(nxt_wr_ptr[2]), 
        .A4(nxt_wr_ptr[30]), .Z(n1883) );
  OR4_X1 U1608 ( .A1(nxt_wr_ptr[31]), .A2(nxt_wr_ptr[32]), .A3(nxt_wr_ptr[33]), 
        .A4(nxt_wr_ptr[34]), .Z(n1884) );
  OR4_X1 U1609 ( .A1(nxt_wr_ptr[35]), .A2(nxt_wr_ptr[36]), .A3(nxt_wr_ptr[37]), 
        .A4(nxt_wr_ptr[38]), .Z(n1885) );
  OR4_X1 U1610 ( .A1(nxt_wr_ptr[13]), .A2(nxt_wr_ptr[14]), .A3(nxt_wr_ptr[15]), 
        .A4(nxt_wr_ptr[16]), .Z(n1879) );
  OR4_X1 U1611 ( .A1(nxt_wr_ptr[17]), .A2(nxt_wr_ptr[18]), .A3(nxt_wr_ptr[19]), 
        .A4(nxt_wr_ptr[1]), .Z(n1880) );
  OR4_X1 U1612 ( .A1(nxt_wr_ptr[20]), .A2(nxt_wr_ptr[21]), .A3(nxt_wr_ptr[22]), 
        .A4(nxt_wr_ptr[23]), .Z(n1881) );
  AND2_X1 U1613 ( .A1(wr), .A2(n1712), .Z(n2216) );
  circ_q_WORD_SZ64_0_DW01_inc_0 add_97 ( .A(nxt_wr_ptr), .SUM({N595, N594, 
        N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, 
        N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, 
        N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, 
        N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, 
        N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, 
        N533, N532}) );
  circ_q_WORD_SZ64_0_DW01_inc_1 add_72 ( .A(nxt_rd_ptr), .SUM({N309, N308, 
        N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, 
        N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, 
        N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, 
        N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, 
        N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, 
        N247, N246}) );
  BUF_X2 U4 ( .I(n950), .Z(n471) );
  BUF_X2 U452 ( .I(n2073), .Z(n484) );
  BUF_X2 U453 ( .I(n2073), .Z(n483) );
  BUF_X2 U454 ( .I(n2073), .Z(n479) );
  BUF_X2 U455 ( .I(n2073), .Z(n480) );
  BUF_X2 U456 ( .I(n2073), .Z(n481) );
  BUF_X2 U457 ( .I(n2073), .Z(n482) );
  BUF_X2 U458 ( .I(n2008), .Z(n477) );
  BUF_X2 U459 ( .I(n2008), .Z(n472) );
  BUF_X2 U460 ( .I(n2008), .Z(n473) );
  BUF_X2 U461 ( .I(n2008), .Z(n474) );
  BUF_X2 U462 ( .I(n2008), .Z(n475) );
  BUF_X2 U463 ( .I(n2008), .Z(n476) );
  BUF_X2 U464 ( .I(n950), .Z(n470) );
  BUF_X2 U465 ( .I(n950), .Z(n469) );
  BUF_X2 U466 ( .I(n950), .Z(n468) );
  BUF_X2 U467 ( .I(n950), .Z(n467) );
  INV_X1 U468 ( .I(n564), .ZN(n532) );
  INV_X1 U469 ( .I(n564), .ZN(n533) );
  INV_X1 U470 ( .I(n564), .ZN(n534) );
  INV_X1 U471 ( .I(n515), .ZN(n524) );
  INV_X1 U472 ( .I(n565), .ZN(n535) );
  INV_X1 U473 ( .I(n565), .ZN(n536) );
  INV_X1 U474 ( .I(n456), .ZN(n950) );
  NAND2_X1 U475 ( .A1(n449), .A2(n2006), .ZN(n2008) );
  BUF_X2 U476 ( .I(n709), .Z(n462) );
  BUF_X2 U477 ( .I(n2367), .Z(n571) );
  BUF_X2 U478 ( .I(n578), .Z(n577) );
  BUF_X2 U479 ( .I(n579), .Z(n573) );
  BUF_X2 U480 ( .I(n579), .Z(n574) );
  BUF_X2 U481 ( .I(n579), .Z(n572) );
  BUF_X2 U482 ( .I(n578), .Z(n575) );
  BUF_X2 U483 ( .I(n578), .Z(n576) );
  INV_X1 U484 ( .I(n449), .ZN(n478) );
  BUF_X2 U485 ( .I(n516), .Z(n515) );
  BUF_X2 U486 ( .I(n2367), .Z(n570) );
  BUF_X2 U487 ( .I(n2367), .Z(n566) );
  BUF_X2 U488 ( .I(n2367), .Z(n567) );
  BUF_X2 U489 ( .I(n2367), .Z(n568) );
  BUF_X2 U490 ( .I(n2367), .Z(n569) );
  INV_X1 U491 ( .I(n493), .ZN(n487) );
  INV_X1 U492 ( .I(n493), .ZN(n489) );
  INV_X1 U493 ( .I(n493), .ZN(n488) );
  BUF_X2 U494 ( .I(n709), .Z(n465) );
  BUF_X2 U495 ( .I(n709), .Z(n464) );
  BUF_X2 U496 ( .I(n709), .Z(n463) );
  BUF_X2 U497 ( .I(n709), .Z(n461) );
  BUF_X2 U498 ( .I(n709), .Z(n460) );
  BUF_X2 U499 ( .I(n709), .Z(n459) );
  BUF_X2 U500 ( .I(n709), .Z(n458) );
  BUF_X2 U501 ( .I(n709), .Z(n457) );
  BUF_X2 U502 ( .I(n516), .Z(n514) );
  BUF_X2 U503 ( .I(n517), .Z(n513) );
  BUF_X2 U504 ( .I(n517), .Z(n512) );
  BUF_X2 U505 ( .I(n517), .Z(n511) );
  BUF_X2 U506 ( .I(n518), .Z(n510) );
  BUF_X2 U507 ( .I(n518), .Z(n509) );
  BUF_X2 U508 ( .I(n518), .Z(n508) );
  BUF_X2 U509 ( .I(n519), .Z(n507) );
  BUF_X2 U510 ( .I(n519), .Z(n506) );
  BUF_X2 U511 ( .I(n519), .Z(n505) );
  BUF_X2 U512 ( .I(n520), .Z(n504) );
  BUF_X2 U513 ( .I(n520), .Z(n503) );
  BUF_X2 U514 ( .I(n520), .Z(n502) );
  BUF_X2 U515 ( .I(n521), .Z(n501) );
  BUF_X2 U516 ( .I(n521), .Z(n500) );
  BUF_X2 U517 ( .I(n521), .Z(n499) );
  BUF_X2 U518 ( .I(n522), .Z(n498) );
  BUF_X2 U519 ( .I(n522), .Z(n497) );
  BUF_X2 U520 ( .I(n522), .Z(n496) );
  BUF_X2 U521 ( .I(n523), .Z(n495) );
  BUF_X2 U522 ( .I(n523), .Z(n494) );
  BUF_X2 U523 ( .I(n709), .Z(n466) );
  INV_X1 U524 ( .I(n492), .ZN(n485) );
  INV_X1 U525 ( .I(n491), .ZN(n486) );
  OAI22_X1 U526 ( .A1(n896), .A2(n462), .B1(n472), .B2(n712), .ZN(n1802) );
  INV_X1 U527 ( .I(N308), .ZN(n712) );
  OAI22_X1 U528 ( .A1(n894), .A2(n462), .B1(n472), .B2(n713), .ZN(n1801) );
  INV_X1 U529 ( .I(N307), .ZN(n713) );
  OAI22_X1 U530 ( .A1(n892), .A2(n462), .B1(n472), .B2(n714), .ZN(n1800) );
  INV_X1 U531 ( .I(N306), .ZN(n714) );
  OAI22_X1 U532 ( .A1(n890), .A2(n462), .B1(n472), .B2(n715), .ZN(n1799) );
  INV_X1 U533 ( .I(N305), .ZN(n715) );
  OAI22_X1 U534 ( .A1(n888), .A2(n461), .B1(n472), .B2(n716), .ZN(n1798) );
  INV_X1 U535 ( .I(N304), .ZN(n716) );
  OAI22_X1 U536 ( .A1(n886), .A2(n461), .B1(n472), .B2(n717), .ZN(n1797) );
  INV_X1 U537 ( .I(N303), .ZN(n717) );
  OAI22_X1 U538 ( .A1(n884), .A2(n461), .B1(n472), .B2(n718), .ZN(n1796) );
  INV_X1 U539 ( .I(N302), .ZN(n718) );
  OAI22_X1 U540 ( .A1(n882), .A2(n461), .B1(n472), .B2(n719), .ZN(n1795) );
  INV_X1 U541 ( .I(N301), .ZN(n719) );
  OAI22_X1 U542 ( .A1(n880), .A2(n461), .B1(n472), .B2(n720), .ZN(n1794) );
  INV_X1 U543 ( .I(N300), .ZN(n720) );
  OAI22_X1 U544 ( .A1(n878), .A2(n461), .B1(n472), .B2(n721), .ZN(n1793) );
  INV_X1 U545 ( .I(N299), .ZN(n721) );
  OAI22_X1 U546 ( .A1(n876), .A2(n461), .B1(n472), .B2(n722), .ZN(n1792) );
  INV_X1 U547 ( .I(N298), .ZN(n722) );
  OAI22_X1 U548 ( .A1(n874), .A2(n461), .B1(n472), .B2(n723), .ZN(n1791) );
  INV_X1 U549 ( .I(N297), .ZN(n723) );
  OAI22_X1 U550 ( .A1(n872), .A2(n461), .B1(n473), .B2(n724), .ZN(n1790) );
  INV_X1 U551 ( .I(N296), .ZN(n724) );
  OAI22_X1 U552 ( .A1(n870), .A2(n461), .B1(n473), .B2(n725), .ZN(n1789) );
  INV_X1 U553 ( .I(N295), .ZN(n725) );
  OAI22_X1 U554 ( .A1(n868), .A2(n461), .B1(n473), .B2(n726), .ZN(n1788) );
  INV_X1 U555 ( .I(N294), .ZN(n726) );
  OAI22_X1 U556 ( .A1(n866), .A2(n461), .B1(n473), .B2(n727), .ZN(n1787) );
  INV_X1 U557 ( .I(N293), .ZN(n727) );
  OAI22_X1 U558 ( .A1(n864), .A2(n460), .B1(n473), .B2(n728), .ZN(n1786) );
  INV_X1 U559 ( .I(N292), .ZN(n728) );
  OAI22_X1 U560 ( .A1(n862), .A2(n460), .B1(n473), .B2(n729), .ZN(n1785) );
  INV_X1 U561 ( .I(N291), .ZN(n729) );
  OAI22_X1 U562 ( .A1(n860), .A2(n460), .B1(n473), .B2(n730), .ZN(n1784) );
  INV_X1 U563 ( .I(N290), .ZN(n730) );
  OAI22_X1 U564 ( .A1(n858), .A2(n460), .B1(n473), .B2(n731), .ZN(n1783) );
  INV_X1 U565 ( .I(N289), .ZN(n731) );
  OAI22_X1 U566 ( .A1(n856), .A2(n460), .B1(n473), .B2(n732), .ZN(n1782) );
  INV_X1 U567 ( .I(N288), .ZN(n732) );
  OAI22_X1 U568 ( .A1(n854), .A2(n460), .B1(n473), .B2(n733), .ZN(n1781) );
  INV_X1 U569 ( .I(N287), .ZN(n733) );
  OAI22_X1 U570 ( .A1(n852), .A2(n460), .B1(n473), .B2(n734), .ZN(n1780) );
  INV_X1 U571 ( .I(N286), .ZN(n734) );
  OAI22_X1 U572 ( .A1(n850), .A2(n460), .B1(n473), .B2(n735), .ZN(n1779) );
  INV_X1 U573 ( .I(N285), .ZN(n735) );
  OAI22_X1 U574 ( .A1(n848), .A2(n460), .B1(n474), .B2(n736), .ZN(n1778) );
  INV_X1 U575 ( .I(N284), .ZN(n736) );
  OAI22_X1 U576 ( .A1(n846), .A2(n460), .B1(n474), .B2(n737), .ZN(n1777) );
  INV_X1 U577 ( .I(N283), .ZN(n737) );
  OAI22_X1 U578 ( .A1(n844), .A2(n460), .B1(n474), .B2(n738), .ZN(n1776) );
  INV_X1 U579 ( .I(N282), .ZN(n738) );
  OAI22_X1 U580 ( .A1(n842), .A2(n460), .B1(n474), .B2(n739), .ZN(n1775) );
  INV_X1 U581 ( .I(N281), .ZN(n739) );
  OAI22_X1 U582 ( .A1(n840), .A2(n459), .B1(n474), .B2(n740), .ZN(n1774) );
  INV_X1 U583 ( .I(N280), .ZN(n740) );
  OAI22_X1 U584 ( .A1(n838), .A2(n459), .B1(n474), .B2(n741), .ZN(n1773) );
  INV_X1 U585 ( .I(N279), .ZN(n741) );
  OAI22_X1 U586 ( .A1(n836), .A2(n459), .B1(n474), .B2(n742), .ZN(n1772) );
  INV_X1 U587 ( .I(N278), .ZN(n742) );
  OAI22_X1 U588 ( .A1(n834), .A2(n459), .B1(n474), .B2(n743), .ZN(n1771) );
  INV_X1 U589 ( .I(N277), .ZN(n743) );
  OAI22_X1 U590 ( .A1(n832), .A2(n459), .B1(n474), .B2(n744), .ZN(n1770) );
  INV_X1 U591 ( .I(N276), .ZN(n744) );
  OAI22_X1 U592 ( .A1(n830), .A2(n459), .B1(n474), .B2(n745), .ZN(n1769) );
  INV_X1 U593 ( .I(N275), .ZN(n745) );
  OAI22_X1 U594 ( .A1(n828), .A2(n459), .B1(n474), .B2(n746), .ZN(n1768) );
  INV_X1 U595 ( .I(N274), .ZN(n746) );
  OAI22_X1 U596 ( .A1(n826), .A2(n459), .B1(n474), .B2(n747), .ZN(n1767) );
  INV_X1 U597 ( .I(N273), .ZN(n747) );
  OAI22_X1 U598 ( .A1(n824), .A2(n459), .B1(n475), .B2(n748), .ZN(n1766) );
  INV_X1 U599 ( .I(N272), .ZN(n748) );
  OAI22_X1 U600 ( .A1(n822), .A2(n459), .B1(n475), .B2(n749), .ZN(n1765) );
  INV_X1 U601 ( .I(N271), .ZN(n749) );
  OAI22_X1 U602 ( .A1(n820), .A2(n459), .B1(n475), .B2(n750), .ZN(n1764) );
  INV_X1 U603 ( .I(N270), .ZN(n750) );
  OAI22_X1 U604 ( .A1(n818), .A2(n459), .B1(n475), .B2(n751), .ZN(n1763) );
  INV_X1 U605 ( .I(N269), .ZN(n751) );
  OAI22_X1 U606 ( .A1(n816), .A2(n458), .B1(n475), .B2(n752), .ZN(n1762) );
  INV_X1 U607 ( .I(N268), .ZN(n752) );
  OAI22_X1 U608 ( .A1(n814), .A2(n458), .B1(n475), .B2(n753), .ZN(n1761) );
  INV_X1 U609 ( .I(N267), .ZN(n753) );
  OAI22_X1 U610 ( .A1(n812), .A2(n458), .B1(n475), .B2(n754), .ZN(n1760) );
  INV_X1 U611 ( .I(N266), .ZN(n754) );
  OAI22_X1 U612 ( .A1(n810), .A2(n458), .B1(n475), .B2(n755), .ZN(n1759) );
  INV_X1 U613 ( .I(N265), .ZN(n755) );
  OAI22_X1 U614 ( .A1(n808), .A2(n458), .B1(n475), .B2(n756), .ZN(n1758) );
  INV_X1 U615 ( .I(N264), .ZN(n756) );
  OAI22_X1 U616 ( .A1(n806), .A2(n458), .B1(n475), .B2(n757), .ZN(n1757) );
  INV_X1 U617 ( .I(N263), .ZN(n757) );
  OAI22_X1 U618 ( .A1(n804), .A2(n458), .B1(n475), .B2(n758), .ZN(n1756) );
  INV_X1 U619 ( .I(N262), .ZN(n758) );
  INV_X1 U620 ( .I(n2127), .ZN(n490) );
  BUF_X2 U621 ( .I(n2116), .Z(n456) );
  NAND2_X1 U622 ( .A1(n490), .A2(n1736), .ZN(n2116) );
  OAI22_X1 U623 ( .A1(n802), .A2(n458), .B1(n475), .B2(n759), .ZN(n1755) );
  INV_X1 U624 ( .I(N261), .ZN(n759) );
  INV_X1 U625 ( .I(n2009), .ZN(n709) );
  AND2_X1 U626 ( .A1(n462), .A2(n1736), .Z(n449) );
  OAI22_X1 U627 ( .A1(n777), .A2(n457), .B1(n477), .B2(n772), .ZN(n1742) );
  INV_X1 U628 ( .I(N248), .ZN(n772) );
  OAI22_X1 U629 ( .A1(n776), .A2(n457), .B1(n477), .B2(n773), .ZN(n1741) );
  INV_X1 U630 ( .I(N247), .ZN(n773) );
  OAI22_X1 U631 ( .A1(n800), .A2(n458), .B1(n476), .B2(n760), .ZN(n1754) );
  INV_X1 U632 ( .I(N260), .ZN(n760) );
  OAI22_X1 U633 ( .A1(n798), .A2(n458), .B1(n476), .B2(n761), .ZN(n1753) );
  INV_X1 U634 ( .I(N259), .ZN(n761) );
  OAI22_X1 U635 ( .A1(n796), .A2(n458), .B1(n476), .B2(n762), .ZN(n1752) );
  INV_X1 U636 ( .I(N258), .ZN(n762) );
  OAI22_X1 U637 ( .A1(n794), .A2(n458), .B1(n476), .B2(n763), .ZN(n1751) );
  INV_X1 U638 ( .I(N257), .ZN(n763) );
  OAI22_X1 U639 ( .A1(n792), .A2(n457), .B1(n476), .B2(n764), .ZN(n1750) );
  INV_X1 U640 ( .I(N256), .ZN(n764) );
  OAI22_X1 U641 ( .A1(n790), .A2(n457), .B1(n476), .B2(n765), .ZN(n1749) );
  INV_X1 U642 ( .I(N255), .ZN(n765) );
  OAI22_X1 U643 ( .A1(n788), .A2(n457), .B1(n476), .B2(n766), .ZN(n1748) );
  INV_X1 U644 ( .I(N254), .ZN(n766) );
  OAI22_X1 U645 ( .A1(n786), .A2(n457), .B1(n476), .B2(n767), .ZN(n1747) );
  INV_X1 U646 ( .I(N253), .ZN(n767) );
  OAI22_X1 U647 ( .A1(n784), .A2(n457), .B1(n476), .B2(n768), .ZN(n1746) );
  INV_X1 U648 ( .I(N252), .ZN(n768) );
  OAI22_X1 U649 ( .A1(n782), .A2(n457), .B1(n476), .B2(n769), .ZN(n1745) );
  INV_X1 U650 ( .I(N251), .ZN(n769) );
  OAI22_X1 U651 ( .A1(n780), .A2(n457), .B1(n476), .B2(n770), .ZN(n1744) );
  INV_X1 U652 ( .I(N250), .ZN(n770) );
  OAI22_X1 U653 ( .A1(n778), .A2(n457), .B1(n476), .B2(n771), .ZN(n1743) );
  INV_X1 U654 ( .I(N249), .ZN(n771) );
  NAND4_X1 U655 ( .A1(n2302), .A2(n2301), .A3(n2300), .A4(n2299), .ZN(n2303)
         );
  NOR4_X1 U656 ( .A1(n2286), .A2(n2285), .A3(n2284), .A4(n2283), .ZN(n2302) );
  NOR4_X1 U657 ( .A1(n2290), .A2(n2289), .A3(n2288), .A4(n2287), .ZN(n2301) );
  BUF_X2 U658 ( .I(n2368), .Z(n579) );
  BUF_X2 U659 ( .I(n2368), .Z(n578) );
  OAI22_X1 U660 ( .A1(n462), .A2(n779), .B1(n778), .B2(n478), .ZN(n1804) );
  OAI22_X1 U661 ( .A1(n464), .A2(n851), .B1(n850), .B2(n478), .ZN(n1840) );
  OAI22_X1 U662 ( .A1(n464), .A2(n849), .B1(n848), .B2(n478), .ZN(n1839) );
  OAI22_X1 U663 ( .A1(n464), .A2(n847), .B1(n846), .B2(n478), .ZN(n1838) );
  OAI22_X1 U664 ( .A1(n464), .A2(n845), .B1(n844), .B2(n478), .ZN(n1837) );
  OAI22_X1 U665 ( .A1(n464), .A2(n843), .B1(n842), .B2(n478), .ZN(n1836) );
  OAI22_X1 U666 ( .A1(n464), .A2(n841), .B1(n840), .B2(n478), .ZN(n1835) );
  OAI22_X1 U667 ( .A1(n464), .A2(n839), .B1(n838), .B2(n478), .ZN(n1834) );
  OAI22_X1 U668 ( .A1(n464), .A2(n837), .B1(n836), .B2(n478), .ZN(n1833) );
  OAI22_X1 U669 ( .A1(n464), .A2(n835), .B1(n834), .B2(n478), .ZN(n1832) );
  OAI22_X1 U670 ( .A1(n464), .A2(n833), .B1(n832), .B2(n478), .ZN(n1831) );
  OAI22_X1 U671 ( .A1(n464), .A2(n831), .B1(n830), .B2(n478), .ZN(n1830) );
  OAI22_X1 U672 ( .A1(n464), .A2(n829), .B1(n828), .B2(n478), .ZN(n1829) );
  OAI22_X1 U673 ( .A1(n464), .A2(n827), .B1(n826), .B2(n478), .ZN(n1828) );
  OAI22_X1 U674 ( .A1(n464), .A2(n825), .B1(n824), .B2(n478), .ZN(n1827) );
  OAI22_X1 U675 ( .A1(n463), .A2(n823), .B1(n822), .B2(n478), .ZN(n1826) );
  OAI22_X1 U676 ( .A1(n463), .A2(n821), .B1(n820), .B2(n478), .ZN(n1825) );
  OAI22_X1 U677 ( .A1(n463), .A2(n819), .B1(n818), .B2(n478), .ZN(n1824) );
  OAI22_X1 U678 ( .A1(n463), .A2(n817), .B1(n816), .B2(n478), .ZN(n1823) );
  OAI22_X1 U679 ( .A1(n463), .A2(n815), .B1(n814), .B2(n478), .ZN(n1822) );
  OAI22_X1 U680 ( .A1(n463), .A2(n813), .B1(n812), .B2(n478), .ZN(n1821) );
  OAI22_X1 U681 ( .A1(n463), .A2(n811), .B1(n810), .B2(n478), .ZN(n1820) );
  OAI22_X1 U682 ( .A1(n463), .A2(n809), .B1(n808), .B2(n478), .ZN(n1819) );
  OAI22_X1 U683 ( .A1(n463), .A2(n807), .B1(n806), .B2(n478), .ZN(n1818) );
  OAI22_X1 U684 ( .A1(n463), .A2(n805), .B1(n804), .B2(n478), .ZN(n1817) );
  OAI22_X1 U685 ( .A1(n463), .A2(n803), .B1(n802), .B2(n478), .ZN(n1816) );
  OAI22_X1 U686 ( .A1(n463), .A2(n801), .B1(n800), .B2(n478), .ZN(n1815) );
  OAI22_X1 U687 ( .A1(n463), .A2(n799), .B1(n798), .B2(n478), .ZN(n1814) );
  OAI22_X1 U688 ( .A1(n463), .A2(n797), .B1(n796), .B2(n478), .ZN(n1813) );
  OAI22_X1 U689 ( .A1(n462), .A2(n795), .B1(n794), .B2(n478), .ZN(n1812) );
  OAI22_X1 U690 ( .A1(n462), .A2(n793), .B1(n792), .B2(n478), .ZN(n1811) );
  OAI22_X1 U691 ( .A1(n462), .A2(n791), .B1(n790), .B2(n478), .ZN(n1810) );
  OAI22_X1 U692 ( .A1(n462), .A2(n789), .B1(n788), .B2(n478), .ZN(n1809) );
  OAI22_X1 U693 ( .A1(n462), .A2(n787), .B1(n786), .B2(n478), .ZN(n1808) );
  OAI22_X1 U694 ( .A1(n462), .A2(n785), .B1(n784), .B2(n478), .ZN(n1807) );
  OAI22_X1 U695 ( .A1(n462), .A2(n783), .B1(n782), .B2(n478), .ZN(n1806) );
  OAI22_X1 U696 ( .A1(n462), .A2(n781), .B1(n780), .B2(n478), .ZN(n1805) );
  OAI22_X1 U697 ( .A1(n466), .A2(n893), .B1(n892), .B2(n478), .ZN(n1861) );
  OAI22_X1 U698 ( .A1(n466), .A2(n887), .B1(n886), .B2(n478), .ZN(n1858) );
  OAI22_X1 U699 ( .A1(n465), .A2(n879), .B1(n878), .B2(n478), .ZN(n1854) );
  OAI22_X1 U700 ( .A1(n465), .A2(n865), .B1(n864), .B2(n478), .ZN(n1847) );
  OAI22_X1 U701 ( .A1(n465), .A2(n857), .B1(n856), .B2(n478), .ZN(n1843) );
  OAI22_X1 U702 ( .A1(n466), .A2(n898), .B1(n775), .B2(n478), .ZN(n1864) );
  OAI22_X1 U703 ( .A1(n466), .A2(n895), .B1(n894), .B2(n478), .ZN(n1862) );
  OAI22_X1 U704 ( .A1(n466), .A2(n889), .B1(n888), .B2(n478), .ZN(n1859) );
  OAI22_X1 U705 ( .A1(n466), .A2(n881), .B1(n880), .B2(n478), .ZN(n1855) );
  OAI22_X1 U706 ( .A1(n465), .A2(n873), .B1(n872), .B2(n478), .ZN(n1851) );
  OAI22_X1 U707 ( .A1(n465), .A2(n867), .B1(n866), .B2(n478), .ZN(n1848) );
  OAI22_X1 U708 ( .A1(n465), .A2(n859), .B1(n858), .B2(n478), .ZN(n1844) );
  OAI22_X1 U709 ( .A1(n466), .A2(n897), .B1(n896), .B2(n478), .ZN(n1863) );
  OAI22_X1 U710 ( .A1(n466), .A2(n891), .B1(n890), .B2(n478), .ZN(n1860) );
  OAI22_X1 U711 ( .A1(n466), .A2(n883), .B1(n882), .B2(n478), .ZN(n1856) );
  OAI22_X1 U712 ( .A1(n465), .A2(n875), .B1(n874), .B2(n478), .ZN(n1852) );
  OAI22_X1 U713 ( .A1(n465), .A2(n869), .B1(n868), .B2(n478), .ZN(n1849) );
  OAI22_X1 U714 ( .A1(n465), .A2(n861), .B1(n860), .B2(n478), .ZN(n1845) );
  OAI22_X1 U715 ( .A1(n465), .A2(n853), .B1(n852), .B2(n478), .ZN(n1841) );
  OAI22_X1 U716 ( .A1(n466), .A2(n885), .B1(n884), .B2(n478), .ZN(n1857) );
  OAI22_X1 U717 ( .A1(n465), .A2(n877), .B1(n876), .B2(n478), .ZN(n1853) );
  OAI22_X1 U718 ( .A1(n465), .A2(n871), .B1(n870), .B2(n478), .ZN(n1850) );
  OAI22_X1 U719 ( .A1(n465), .A2(n863), .B1(n862), .B2(n478), .ZN(n1846) );
  OAI22_X1 U720 ( .A1(n465), .A2(n855), .B1(n854), .B2(n478), .ZN(n1842) );
  BUF_X2 U721 ( .I(n2281), .Z(n531) );
  BUF_X2 U722 ( .I(n2213), .Z(n516) );
  INV_X1 U723 ( .I(n2127), .ZN(n493) );
  NOR4_X1 U724 ( .A1(n2298), .A2(n2297), .A3(n2296), .A4(n2295), .ZN(n2299) );
  NAND4_X1 U725 ( .A1(n785), .A2(n787), .A3(n789), .A4(n791), .ZN(n2298) );
  NAND4_X1 U726 ( .A1(n893), .A2(n895), .A3(n897), .A4(n898), .ZN(n2297) );
  NAND4_X1 U727 ( .A1(n887), .A2(n889), .A3(n891), .A4(n783), .ZN(n2296) );
  NAND4_X1 U728 ( .A1(n879), .A2(n881), .A3(n883), .A4(n885), .ZN(n2295) );
  NOR4_X1 U729 ( .A1(n2294), .A2(n2293), .A3(n2292), .A4(n2291), .ZN(n2300) );
  NAND4_X1 U730 ( .A1(n781), .A2(n873), .A3(n875), .A4(n877), .ZN(n2294) );
  NAND4_X1 U731 ( .A1(n865), .A2(n867), .A3(n869), .A4(n871), .ZN(n2293) );
  NAND4_X1 U732 ( .A1(n857), .A2(n859), .A3(n861), .A4(n863), .ZN(n2292) );
  NAND4_X1 U733 ( .A1(n851), .A2(n779), .A3(n853), .A4(n855), .ZN(n2291) );
  NAND4_X1 U734 ( .A1(n819), .A2(n821), .A3(n823), .A4(n825), .ZN(n2287) );
  NAND4_X1 U735 ( .A1(n827), .A2(n829), .A3(n831), .A4(n833), .ZN(n2288) );
  NAND4_X1 U736 ( .A1(n795), .A2(n797), .A3(n799), .A4(n801), .ZN(n2284) );
  NAND4_X1 U737 ( .A1(n835), .A2(n837), .A3(n839), .A4(n841), .ZN(n2289) );
  NAND4_X1 U738 ( .A1(n803), .A2(n805), .A3(n807), .A4(n809), .ZN(n2285) );
  NAND4_X1 U739 ( .A1(n843), .A2(n845), .A3(n847), .A4(n849), .ZN(n2290) );
  OAI22_X1 U740 ( .A1(n492), .A2(n1712), .B1(n456), .B2(n2011), .ZN(n1865) );
  OAI22_X1 U741 ( .A1(n490), .A2(n1733), .B1(n456), .B2(n1732), .ZN(n1876) );
  OAI22_X1 U742 ( .A1(n493), .A2(n1735), .B1(n456), .B2(n1734), .ZN(n1877) );
  OAI22_X1 U743 ( .A1(n492), .A2(n1731), .B1(n456), .B2(n1730), .ZN(n1875) );
  OAI22_X1 U744 ( .A1(n491), .A2(n1729), .B1(n456), .B2(n1728), .ZN(n1874) );
  OAI22_X1 U745 ( .A1(n491), .A2(n1727), .B1(n456), .B2(n1726), .ZN(n1873) );
  OAI22_X1 U746 ( .A1(n491), .A2(n1725), .B1(n456), .B2(n1724), .ZN(n1872) );
  OAI22_X1 U747 ( .A1(n492), .A2(n1723), .B1(n456), .B2(n1722), .ZN(n1871) );
  OAI22_X1 U748 ( .A1(n493), .A2(n1721), .B1(n456), .B2(n1720), .ZN(n1870) );
  OAI22_X1 U749 ( .A1(n492), .A2(n1719), .B1(n456), .B2(n1718), .ZN(n1869) );
  OAI22_X1 U750 ( .A1(n492), .A2(n1717), .B1(n456), .B2(n1716), .ZN(n1868) );
  OAI22_X1 U751 ( .A1(n491), .A2(n1715), .B1(n456), .B2(n1714), .ZN(n1867) );
  BUF_X2 U752 ( .I(n2213), .Z(n517) );
  BUF_X2 U753 ( .I(n2213), .Z(n518) );
  BUF_X2 U754 ( .I(n2213), .Z(n519) );
  BUF_X2 U755 ( .I(n2213), .Z(n520) );
  BUF_X2 U756 ( .I(n2213), .Z(n521) );
  BUF_X2 U757 ( .I(n2213), .Z(n522) );
  BUF_X2 U758 ( .I(n2213), .Z(n523) );
  NAND4_X1 U759 ( .A1(n811), .A2(n813), .A3(n815), .A4(n817), .ZN(n2286) );
  INV_X1 U760 ( .I(n2127), .ZN(n491) );
  INV_X1 U761 ( .I(n2127), .ZN(n492) );
  BUF_X2 U762 ( .I(n2281), .Z(n530) );
  BUF_X2 U763 ( .I(n2281), .Z(n529) );
  BUF_X2 U764 ( .I(n2281), .Z(n528) );
  BUF_X2 U765 ( .I(n2281), .Z(n527) );
  BUF_X2 U766 ( .I(n2281), .Z(n526) );
  BUF_X2 U767 ( .I(n2281), .Z(n525) );
  NAND4_X1 U768 ( .A1(n1723), .A2(n1725), .A3(n1727), .A4(n1729), .ZN(n2143)
         );
  NAND4_X1 U769 ( .A1(n1715), .A2(n1731), .A3(n1733), .A4(n1735), .ZN(n2144)
         );
  NAND4_X1 U770 ( .A1(n1897), .A2(n1896), .A3(n1895), .A4(n1894), .ZN(n1899)
         );
  NOR4_X1 U771 ( .A1(n1881), .A2(n1880), .A3(n1879), .A4(n1878), .ZN(n1897) );
  NOR4_X1 U772 ( .A1(n1885), .A2(n1884), .A3(n1883), .A4(n1882), .ZN(n1896) );
  NOR4_X1 U773 ( .A1(n1889), .A2(n1888), .A3(n1887), .A4(n1886), .ZN(n1895) );
  NAND4_X1 U774 ( .A1(n1722), .A2(n1724), .A3(n1726), .A4(n1728), .ZN(n1888)
         );
  NAND4_X1 U775 ( .A1(n1714), .A2(n1730), .A3(n1732), .A4(n1734), .ZN(n1889)
         );
  OAI21_X1 U776 ( .A1(n2009), .A2(n1985), .B(n710), .ZN(n1738) );
  NAND4_X1 U777 ( .A1(n2005), .A2(n2004), .A3(n2003), .A4(n2002), .ZN(n2006)
         );
  NOR4_X1 U778 ( .A1(n1989), .A2(n1988), .A3(n1987), .A4(n1986), .ZN(n2005) );
  NOR4_X1 U779 ( .A1(n1993), .A2(n1992), .A3(n1991), .A4(n1990), .ZN(n2004) );
  NOR4_X1 U780 ( .A1(n1997), .A2(n1996), .A3(n1995), .A4(n1994), .ZN(n2003) );
  NOR4_X1 U781 ( .A1(n2001), .A2(n2000), .A3(n1999), .A4(n1998), .ZN(n2002) );
  NAND4_X1 U782 ( .A1(n784), .A2(n786), .A3(n788), .A4(n790), .ZN(n2001) );
  NAND4_X1 U783 ( .A1(n886), .A2(n888), .A3(n890), .A4(n782), .ZN(n1999) );
  NAND4_X1 U784 ( .A1(n878), .A2(n880), .A3(n882), .A4(n884), .ZN(n1998) );
  NAND4_X1 U785 ( .A1(n850), .A2(n778), .A3(n852), .A4(n854), .ZN(n1994) );
  NAND4_X1 U786 ( .A1(n892), .A2(n894), .A3(n896), .A4(n775), .ZN(n2000) );
  NAND4_X1 U787 ( .A1(n820), .A2(n822), .A3(n824), .A4(n826), .ZN(n1990) );
  NAND4_X1 U788 ( .A1(n856), .A2(n858), .A3(n860), .A4(n862), .ZN(n1995) );
  NAND4_X1 U789 ( .A1(n828), .A2(n830), .A3(n777), .A4(n832), .ZN(n1991) );
  NAND4_X1 U790 ( .A1(n864), .A2(n866), .A3(n868), .A4(n870), .ZN(n1996) );
  NAND4_X1 U791 ( .A1(n834), .A2(n836), .A3(n838), .A4(n840), .ZN(n1992) );
  NAND4_X1 U792 ( .A1(n798), .A2(n800), .A3(n802), .A4(n804), .ZN(n1987) );
  NAND4_X1 U793 ( .A1(n806), .A2(n808), .A3(n810), .A4(n776), .ZN(n1988) );
  NAND4_X1 U794 ( .A1(n780), .A2(n872), .A3(n874), .A4(n876), .ZN(n1997) );
  NAND4_X1 U795 ( .A1(n842), .A2(n844), .A3(n846), .A4(n848), .ZN(n1993) );
  NAND4_X1 U796 ( .A1(n812), .A2(n814), .A3(n816), .A4(n818), .ZN(n1989) );
  NAND4_X1 U797 ( .A1(n1984), .A2(n1983), .A3(n1982), .A4(n1981), .ZN(n2011)
         );
  NOR4_X1 U798 ( .A1(n1940), .A2(n1939), .A3(n1938), .A4(n1937), .ZN(n1983) );
  NOR4_X1 U799 ( .A1(n1960), .A2(n1959), .A3(n1958), .A4(n1957), .ZN(n1982) );
  NOR4_X1 U800 ( .A1(n1980), .A2(n1979), .A3(n1978), .A4(n1977), .ZN(n1981) );
  NOR4_X1 U801 ( .A1(n1920), .A2(n1919), .A3(n1918), .A4(n1917), .ZN(n1984) );
  NAND4_X1 U802 ( .A1(n1904), .A2(n1903), .A3(n1902), .A4(n1901), .ZN(n1920)
         );
  NAND4_X1 U803 ( .A1(n1908), .A2(n1907), .A3(n1906), .A4(n1905), .ZN(n1919)
         );
  NAND4_X1 U804 ( .A1(n1912), .A2(n1911), .A3(n1910), .A4(n1909), .ZN(n1918)
         );
  INV_X1 U805 ( .I(n1900), .ZN(n580) );
  AOI22_X1 U806 ( .A1(N595), .A2(n484), .B1(n487), .B2(nxt_wr_ptr[63]), .ZN(
        n1900) );
  OAI22_X1 U807 ( .A1(n775), .A2(n457), .B1(n477), .B2(n711), .ZN(n1739) );
  INV_X1 U808 ( .I(N309), .ZN(n711) );
  INV_X1 U809 ( .I(n2074), .ZN(n581) );
  AOI22_X1 U810 ( .A1(N594), .A2(n479), .B1(nxt_wr_ptr[62]), .B2(n489), .ZN(
        n2074) );
  INV_X1 U811 ( .I(n2072), .ZN(n582) );
  AOI22_X1 U812 ( .A1(N593), .A2(n479), .B1(nxt_wr_ptr[61]), .B2(n488), .ZN(
        n2072) );
  INV_X1 U813 ( .I(n2071), .ZN(n583) );
  AOI22_X1 U814 ( .A1(N592), .A2(n479), .B1(nxt_wr_ptr[60]), .B2(n487), .ZN(
        n2071) );
  INV_X1 U815 ( .I(n2070), .ZN(n584) );
  AOI22_X1 U816 ( .A1(N591), .A2(n479), .B1(nxt_wr_ptr[59]), .B2(n486), .ZN(
        n2070) );
  INV_X1 U817 ( .I(n2069), .ZN(n585) );
  AOI22_X1 U818 ( .A1(N590), .A2(n479), .B1(nxt_wr_ptr[58]), .B2(n487), .ZN(
        n2069) );
  INV_X1 U819 ( .I(n2068), .ZN(n586) );
  AOI22_X1 U820 ( .A1(N589), .A2(n479), .B1(nxt_wr_ptr[57]), .B2(n485), .ZN(
        n2068) );
  INV_X1 U821 ( .I(n2067), .ZN(n587) );
  AOI22_X1 U822 ( .A1(N588), .A2(n479), .B1(nxt_wr_ptr[56]), .B2(n487), .ZN(
        n2067) );
  INV_X1 U823 ( .I(n2066), .ZN(n588) );
  AOI22_X1 U824 ( .A1(N587), .A2(n479), .B1(nxt_wr_ptr[55]), .B2(n489), .ZN(
        n2066) );
  INV_X1 U825 ( .I(n2065), .ZN(n589) );
  AOI22_X1 U826 ( .A1(N586), .A2(n479), .B1(nxt_wr_ptr[54]), .B2(n488), .ZN(
        n2065) );
  INV_X1 U827 ( .I(n2064), .ZN(n590) );
  AOI22_X1 U828 ( .A1(N585), .A2(n479), .B1(nxt_wr_ptr[53]), .B2(n485), .ZN(
        n2064) );
  INV_X1 U829 ( .I(n2063), .ZN(n591) );
  AOI22_X1 U830 ( .A1(N584), .A2(n479), .B1(nxt_wr_ptr[52]), .B2(n486), .ZN(
        n2063) );
  INV_X1 U831 ( .I(n2062), .ZN(n592) );
  AOI22_X1 U832 ( .A1(N583), .A2(n479), .B1(nxt_wr_ptr[51]), .B2(n486), .ZN(
        n2062) );
  INV_X1 U833 ( .I(n2061), .ZN(n593) );
  AOI22_X1 U834 ( .A1(N582), .A2(n480), .B1(nxt_wr_ptr[50]), .B2(n486), .ZN(
        n2061) );
  INV_X1 U835 ( .I(n2060), .ZN(n594) );
  AOI22_X1 U836 ( .A1(N581), .A2(n480), .B1(nxt_wr_ptr[49]), .B2(n489), .ZN(
        n2060) );
  INV_X1 U837 ( .I(n2059), .ZN(n595) );
  AOI22_X1 U838 ( .A1(N580), .A2(n480), .B1(nxt_wr_ptr[48]), .B2(n488), .ZN(
        n2059) );
  INV_X1 U839 ( .I(n2058), .ZN(n596) );
  AOI22_X1 U840 ( .A1(N579), .A2(n480), .B1(nxt_wr_ptr[47]), .B2(n486), .ZN(
        n2058) );
  INV_X1 U841 ( .I(n2057), .ZN(n597) );
  AOI22_X1 U842 ( .A1(N578), .A2(n480), .B1(nxt_wr_ptr[46]), .B2(n485), .ZN(
        n2057) );
  INV_X1 U843 ( .I(n2056), .ZN(n598) );
  AOI22_X1 U844 ( .A1(N577), .A2(n480), .B1(nxt_wr_ptr[45]), .B2(n489), .ZN(
        n2056) );
  INV_X1 U845 ( .I(n2055), .ZN(n599) );
  AOI22_X1 U846 ( .A1(N576), .A2(n480), .B1(nxt_wr_ptr[44]), .B2(n488), .ZN(
        n2055) );
  INV_X1 U847 ( .I(n2054), .ZN(n600) );
  AOI22_X1 U848 ( .A1(N575), .A2(n480), .B1(nxt_wr_ptr[43]), .B2(n487), .ZN(
        n2054) );
  INV_X1 U849 ( .I(n2053), .ZN(n601) );
  AOI22_X1 U850 ( .A1(N574), .A2(n480), .B1(nxt_wr_ptr[42]), .B2(n486), .ZN(
        n2053) );
  INV_X1 U851 ( .I(n2052), .ZN(n602) );
  AOI22_X1 U852 ( .A1(N573), .A2(n480), .B1(nxt_wr_ptr[41]), .B2(n485), .ZN(
        n2052) );
  INV_X1 U853 ( .I(n2051), .ZN(n603) );
  AOI22_X1 U854 ( .A1(N572), .A2(n480), .B1(nxt_wr_ptr[40]), .B2(n489), .ZN(
        n2051) );
  INV_X1 U855 ( .I(n2050), .ZN(n604) );
  AOI22_X1 U856 ( .A1(N571), .A2(n480), .B1(nxt_wr_ptr[39]), .B2(n488), .ZN(
        n2050) );
  INV_X1 U857 ( .I(n2049), .ZN(n605) );
  AOI22_X1 U858 ( .A1(N570), .A2(n481), .B1(nxt_wr_ptr[38]), .B2(n485), .ZN(
        n2049) );
  INV_X1 U859 ( .I(n2048), .ZN(n606) );
  AOI22_X1 U860 ( .A1(N569), .A2(n481), .B1(nxt_wr_ptr[37]), .B2(n485), .ZN(
        n2048) );
  INV_X1 U861 ( .I(n2047), .ZN(n607) );
  AOI22_X1 U862 ( .A1(N568), .A2(n481), .B1(nxt_wr_ptr[36]), .B2(n485), .ZN(
        n2047) );
  INV_X1 U863 ( .I(n2046), .ZN(n608) );
  AOI22_X1 U864 ( .A1(N567), .A2(n481), .B1(nxt_wr_ptr[35]), .B2(n485), .ZN(
        n2046) );
  INV_X1 U865 ( .I(n2045), .ZN(n609) );
  AOI22_X1 U866 ( .A1(N566), .A2(n481), .B1(nxt_wr_ptr[34]), .B2(n485), .ZN(
        n2045) );
  INV_X1 U867 ( .I(n2044), .ZN(n610) );
  AOI22_X1 U868 ( .A1(N565), .A2(n481), .B1(nxt_wr_ptr[33]), .B2(n485), .ZN(
        n2044) );
  INV_X1 U869 ( .I(n2043), .ZN(n611) );
  AOI22_X1 U870 ( .A1(N564), .A2(n481), .B1(nxt_wr_ptr[32]), .B2(n485), .ZN(
        n2043) );
  INV_X1 U871 ( .I(n2042), .ZN(n612) );
  AOI22_X1 U872 ( .A1(N563), .A2(n481), .B1(nxt_wr_ptr[31]), .B2(n485), .ZN(
        n2042) );
  INV_X1 U873 ( .I(n2041), .ZN(n613) );
  AOI22_X1 U874 ( .A1(N562), .A2(n481), .B1(nxt_wr_ptr[30]), .B2(n485), .ZN(
        n2041) );
  INV_X1 U875 ( .I(n2040), .ZN(n614) );
  AOI22_X1 U876 ( .A1(N561), .A2(n481), .B1(nxt_wr_ptr[29]), .B2(n485), .ZN(
        n2040) );
  INV_X1 U877 ( .I(n2039), .ZN(n615) );
  AOI22_X1 U878 ( .A1(N560), .A2(n481), .B1(nxt_wr_ptr[28]), .B2(n485), .ZN(
        n2039) );
  INV_X1 U879 ( .I(n2038), .ZN(n616) );
  AOI22_X1 U880 ( .A1(N559), .A2(n481), .B1(nxt_wr_ptr[27]), .B2(n485), .ZN(
        n2038) );
  INV_X1 U881 ( .I(n2037), .ZN(n617) );
  AOI22_X1 U882 ( .A1(N558), .A2(n482), .B1(nxt_wr_ptr[26]), .B2(n486), .ZN(
        n2037) );
  INV_X1 U883 ( .I(n2036), .ZN(n618) );
  AOI22_X1 U884 ( .A1(N557), .A2(n482), .B1(nxt_wr_ptr[25]), .B2(n486), .ZN(
        n2036) );
  INV_X1 U885 ( .I(n2035), .ZN(n619) );
  AOI22_X1 U886 ( .A1(N556), .A2(n482), .B1(nxt_wr_ptr[24]), .B2(n486), .ZN(
        n2035) );
  INV_X1 U887 ( .I(n2034), .ZN(n620) );
  AOI22_X1 U888 ( .A1(N555), .A2(n482), .B1(nxt_wr_ptr[23]), .B2(n486), .ZN(
        n2034) );
  INV_X1 U889 ( .I(n2033), .ZN(n621) );
  AOI22_X1 U890 ( .A1(N554), .A2(n482), .B1(nxt_wr_ptr[22]), .B2(n486), .ZN(
        n2033) );
  INV_X1 U891 ( .I(n2032), .ZN(n622) );
  AOI22_X1 U892 ( .A1(N553), .A2(n482), .B1(nxt_wr_ptr[21]), .B2(n486), .ZN(
        n2032) );
  INV_X1 U893 ( .I(n2031), .ZN(n623) );
  AOI22_X1 U894 ( .A1(N552), .A2(n482), .B1(nxt_wr_ptr[20]), .B2(n486), .ZN(
        n2031) );
  INV_X1 U895 ( .I(n2030), .ZN(n624) );
  AOI22_X1 U896 ( .A1(N551), .A2(n482), .B1(nxt_wr_ptr[19]), .B2(n486), .ZN(
        n2030) );
  INV_X1 U897 ( .I(n2029), .ZN(n625) );
  AOI22_X1 U898 ( .A1(N550), .A2(n482), .B1(nxt_wr_ptr[18]), .B2(n486), .ZN(
        n2029) );
  INV_X1 U899 ( .I(n2028), .ZN(n626) );
  AOI22_X1 U900 ( .A1(N549), .A2(n482), .B1(nxt_wr_ptr[17]), .B2(n486), .ZN(
        n2028) );
  INV_X1 U901 ( .I(n2027), .ZN(n627) );
  AOI22_X1 U902 ( .A1(N548), .A2(n482), .B1(nxt_wr_ptr[16]), .B2(n486), .ZN(
        n2027) );
  NOR2_X1 U903 ( .A1(rst), .A2(n2216), .ZN(n2127) );
  INV_X1 U904 ( .I(n2024), .ZN(n630) );
  AOI22_X1 U905 ( .A1(N545), .A2(n483), .B1(nxt_wr_ptr[13]), .B2(n487), .ZN(
        n2024) );
  INV_X1 U906 ( .I(n2017), .ZN(n637) );
  AOI22_X1 U907 ( .A1(N538), .A2(n483), .B1(nxt_wr_ptr[6]), .B2(n486), .ZN(
        n2017) );
  INV_X1 U908 ( .I(n2025), .ZN(n629) );
  AOI22_X1 U909 ( .A1(N546), .A2(n483), .B1(nxt_wr_ptr[14]), .B2(n489), .ZN(
        n2025) );
  INV_X1 U910 ( .I(n2018), .ZN(n636) );
  AOI22_X1 U911 ( .A1(N539), .A2(n483), .B1(nxt_wr_ptr[7]), .B2(n488), .ZN(
        n2018) );
  INV_X1 U912 ( .I(n2014), .ZN(n640) );
  AOI22_X1 U913 ( .A1(N535), .A2(n483), .B1(nxt_wr_ptr[3]), .B2(n485), .ZN(
        n2014) );
  INV_X1 U914 ( .I(n2026), .ZN(n628) );
  AOI22_X1 U915 ( .A1(N547), .A2(n482), .B1(nxt_wr_ptr[15]), .B2(n486), .ZN(
        n2026) );
  INV_X1 U916 ( .I(n2019), .ZN(n635) );
  AOI22_X1 U917 ( .A1(N540), .A2(n483), .B1(nxt_wr_ptr[8]), .B2(n487), .ZN(
        n2019) );
  INV_X1 U918 ( .I(n2013), .ZN(n641) );
  AOI22_X1 U919 ( .A1(N534), .A2(n484), .B1(nxt_wr_ptr[2]), .B2(n487), .ZN(
        n2013) );
  INV_X1 U920 ( .I(n2020), .ZN(n634) );
  AOI22_X1 U921 ( .A1(N541), .A2(n483), .B1(nxt_wr_ptr[9]), .B2(n486), .ZN(
        n2020) );
  INV_X1 U922 ( .I(n2016), .ZN(n638) );
  AOI22_X1 U923 ( .A1(N537), .A2(n483), .B1(nxt_wr_ptr[5]), .B2(n489), .ZN(
        n2016) );
  INV_X1 U924 ( .I(n2012), .ZN(n642) );
  AOI22_X1 U925 ( .A1(N533), .A2(n484), .B1(nxt_wr_ptr[1]), .B2(n487), .ZN(
        n2012) );
  INV_X1 U926 ( .I(n2023), .ZN(n631) );
  AOI22_X1 U927 ( .A1(N544), .A2(n483), .B1(nxt_wr_ptr[12]), .B2(n488), .ZN(
        n2023) );
  INV_X1 U928 ( .I(n2022), .ZN(n632) );
  AOI22_X1 U929 ( .A1(N543), .A2(n483), .B1(nxt_wr_ptr[11]), .B2(n485), .ZN(
        n2022) );
  INV_X1 U930 ( .I(n2021), .ZN(n633) );
  AOI22_X1 U931 ( .A1(N542), .A2(n483), .B1(nxt_wr_ptr[10]), .B2(n485), .ZN(
        n2021) );
  INV_X1 U932 ( .I(n2015), .ZN(n639) );
  AOI22_X1 U933 ( .A1(N536), .A2(n483), .B1(nxt_wr_ptr[4]), .B2(n487), .ZN(
        n2015) );
  AOI21_X1 U934 ( .A1(n710), .A2(rd), .B(rst), .ZN(n2009) );
  INV_X1 U935 ( .I(rst), .ZN(n1736) );
  NOR2_X1 U936 ( .A1(n571), .A2(rst), .ZN(n2368) );
  INV_X1 U937 ( .I(n2335), .ZN(n676) );
  AOI22_X1 U938 ( .A1(N214), .A2(n574), .B1(data_out[32]), .B2(n568), .ZN(
        n2335) );
  INV_X1 U939 ( .I(n2334), .ZN(n675) );
  AOI22_X1 U940 ( .A1(N215), .A2(n574), .B1(data_out[33]), .B2(n568), .ZN(
        n2334) );
  INV_X1 U941 ( .I(n2332), .ZN(n673) );
  AOI22_X1 U942 ( .A1(N217), .A2(n574), .B1(data_out[35]), .B2(n568), .ZN(
        n2332) );
  INV_X1 U943 ( .I(n2333), .ZN(n674) );
  AOI22_X1 U944 ( .A1(N216), .A2(n574), .B1(data_out[34]), .B2(n568), .ZN(
        n2333) );
  INV_X1 U945 ( .I(n2307), .ZN(n648) );
  AOI22_X1 U946 ( .A1(N242), .A2(n577), .B1(data_out[60]), .B2(n571), .ZN(
        n2307) );
  INV_X1 U947 ( .I(n2306), .ZN(n647) );
  AOI22_X1 U948 ( .A1(N243), .A2(n577), .B1(data_out[61]), .B2(n571), .ZN(
        n2306) );
  INV_X1 U949 ( .I(n2305), .ZN(n646) );
  AOI22_X1 U950 ( .A1(N244), .A2(n577), .B1(data_out[62]), .B2(n571), .ZN(
        n2305) );
  INV_X1 U951 ( .I(n2304), .ZN(n645) );
  AOI22_X1 U952 ( .A1(N245), .A2(n577), .B1(data_out[63]), .B2(n571), .ZN(
        n2304) );
  INV_X1 U953 ( .I(n2369), .ZN(n708) );
  AOI22_X1 U954 ( .A1(N182), .A2(n572), .B1(data_out[0]), .B2(n566), .ZN(n2369) );
  INV_X1 U955 ( .I(n2366), .ZN(n707) );
  AOI22_X1 U956 ( .A1(N183), .A2(n572), .B1(data_out[1]), .B2(n566), .ZN(n2366) );
  INV_X1 U957 ( .I(n2365), .ZN(n706) );
  AOI22_X1 U958 ( .A1(N184), .A2(n572), .B1(data_out[2]), .B2(n566), .ZN(n2365) );
  INV_X1 U959 ( .I(n2364), .ZN(n705) );
  AOI22_X1 U960 ( .A1(N185), .A2(n572), .B1(data_out[3]), .B2(n566), .ZN(n2364) );
  INV_X1 U961 ( .I(n2363), .ZN(n704) );
  AOI22_X1 U962 ( .A1(N186), .A2(n572), .B1(data_out[4]), .B2(n566), .ZN(n2363) );
  INV_X1 U963 ( .I(n2362), .ZN(n703) );
  AOI22_X1 U964 ( .A1(N187), .A2(n572), .B1(data_out[5]), .B2(n566), .ZN(n2362) );
  INV_X1 U965 ( .I(n2361), .ZN(n702) );
  AOI22_X1 U966 ( .A1(N188), .A2(n572), .B1(data_out[6]), .B2(n566), .ZN(n2361) );
  INV_X1 U967 ( .I(n2360), .ZN(n701) );
  AOI22_X1 U968 ( .A1(N189), .A2(n572), .B1(data_out[7]), .B2(n566), .ZN(n2360) );
  INV_X1 U969 ( .I(n2359), .ZN(n700) );
  AOI22_X1 U970 ( .A1(N190), .A2(n572), .B1(data_out[8]), .B2(n566), .ZN(n2359) );
  INV_X1 U971 ( .I(n2358), .ZN(n699) );
  AOI22_X1 U972 ( .A1(N191), .A2(n572), .B1(data_out[9]), .B2(n566), .ZN(n2358) );
  INV_X1 U973 ( .I(n2357), .ZN(n698) );
  AOI22_X1 U974 ( .A1(N192), .A2(n572), .B1(data_out[10]), .B2(n566), .ZN(
        n2357) );
  INV_X1 U975 ( .I(n2356), .ZN(n697) );
  AOI22_X1 U976 ( .A1(N193), .A2(n572), .B1(data_out[11]), .B2(n566), .ZN(
        n2356) );
  INV_X1 U977 ( .I(n2355), .ZN(n696) );
  AOI22_X1 U978 ( .A1(N194), .A2(n573), .B1(data_out[12]), .B2(n567), .ZN(
        n2355) );
  INV_X1 U979 ( .I(n2354), .ZN(n695) );
  AOI22_X1 U980 ( .A1(N195), .A2(n573), .B1(data_out[13]), .B2(n567), .ZN(
        n2354) );
  INV_X1 U981 ( .I(n2353), .ZN(n694) );
  AOI22_X1 U982 ( .A1(N196), .A2(n573), .B1(data_out[14]), .B2(n567), .ZN(
        n2353) );
  INV_X1 U983 ( .I(n2352), .ZN(n693) );
  AOI22_X1 U984 ( .A1(N197), .A2(n573), .B1(data_out[15]), .B2(n567), .ZN(
        n2352) );
  INV_X1 U985 ( .I(n2351), .ZN(n692) );
  AOI22_X1 U986 ( .A1(N198), .A2(n573), .B1(data_out[16]), .B2(n567), .ZN(
        n2351) );
  INV_X1 U987 ( .I(n2350), .ZN(n691) );
  AOI22_X1 U988 ( .A1(N199), .A2(n573), .B1(data_out[17]), .B2(n567), .ZN(
        n2350) );
  INV_X1 U989 ( .I(n2349), .ZN(n690) );
  AOI22_X1 U990 ( .A1(N200), .A2(n573), .B1(data_out[18]), .B2(n567), .ZN(
        n2349) );
  INV_X1 U991 ( .I(n2348), .ZN(n689) );
  AOI22_X1 U992 ( .A1(N201), .A2(n573), .B1(data_out[19]), .B2(n567), .ZN(
        n2348) );
  INV_X1 U993 ( .I(n2347), .ZN(n688) );
  AOI22_X1 U994 ( .A1(N202), .A2(n573), .B1(data_out[20]), .B2(n567), .ZN(
        n2347) );
  INV_X1 U995 ( .I(n2346), .ZN(n687) );
  AOI22_X1 U996 ( .A1(N203), .A2(n573), .B1(data_out[21]), .B2(n567), .ZN(
        n2346) );
  INV_X1 U997 ( .I(n2345), .ZN(n686) );
  AOI22_X1 U998 ( .A1(N204), .A2(n573), .B1(data_out[22]), .B2(n567), .ZN(
        n2345) );
  INV_X1 U999 ( .I(n2344), .ZN(n685) );
  AOI22_X1 U1000 ( .A1(N205), .A2(n573), .B1(data_out[23]), .B2(n567), .ZN(
        n2344) );
  INV_X1 U1001 ( .I(n2343), .ZN(n684) );
  AOI22_X1 U1002 ( .A1(N206), .A2(n574), .B1(data_out[24]), .B2(n568), .ZN(
        n2343) );
  INV_X1 U1003 ( .I(n2342), .ZN(n683) );
  AOI22_X1 U1004 ( .A1(N207), .A2(n574), .B1(data_out[25]), .B2(n568), .ZN(
        n2342) );
  INV_X1 U1005 ( .I(n2341), .ZN(n682) );
  AOI22_X1 U1006 ( .A1(N208), .A2(n574), .B1(data_out[26]), .B2(n568), .ZN(
        n2341) );
  INV_X1 U1007 ( .I(n2340), .ZN(n681) );
  AOI22_X1 U1008 ( .A1(N209), .A2(n574), .B1(data_out[27]), .B2(n568), .ZN(
        n2340) );
  INV_X1 U1009 ( .I(n2339), .ZN(n680) );
  AOI22_X1 U1010 ( .A1(N210), .A2(n574), .B1(data_out[28]), .B2(n568), .ZN(
        n2339) );
  INV_X1 U1011 ( .I(n2338), .ZN(n679) );
  AOI22_X1 U1012 ( .A1(N211), .A2(n574), .B1(data_out[29]), .B2(n568), .ZN(
        n2338) );
  INV_X1 U1013 ( .I(n2337), .ZN(n678) );
  AOI22_X1 U1014 ( .A1(N212), .A2(n574), .B1(data_out[30]), .B2(n568), .ZN(
        n2337) );
  INV_X1 U1015 ( .I(n2336), .ZN(n677) );
  AOI22_X1 U1016 ( .A1(N213), .A2(n574), .B1(data_out[31]), .B2(n568), .ZN(
        n2336) );
  INV_X1 U1017 ( .I(n2330), .ZN(n671) );
  AOI22_X1 U1018 ( .A1(N219), .A2(n575), .B1(data_out[37]), .B2(n569), .ZN(
        n2330) );
  INV_X1 U1019 ( .I(n2328), .ZN(n669) );
  AOI22_X1 U1020 ( .A1(N221), .A2(n575), .B1(data_out[39]), .B2(n569), .ZN(
        n2328) );
  INV_X1 U1021 ( .I(n2327), .ZN(n668) );
  AOI22_X1 U1022 ( .A1(N222), .A2(n575), .B1(data_out[40]), .B2(n569), .ZN(
        n2327) );
  INV_X1 U1023 ( .I(n2326), .ZN(n667) );
  AOI22_X1 U1024 ( .A1(N223), .A2(n575), .B1(data_out[41]), .B2(n569), .ZN(
        n2326) );
  INV_X1 U1025 ( .I(n2324), .ZN(n665) );
  AOI22_X1 U1026 ( .A1(N225), .A2(n575), .B1(data_out[43]), .B2(n569), .ZN(
        n2324) );
  INV_X1 U1027 ( .I(n2322), .ZN(n663) );
  AOI22_X1 U1028 ( .A1(N227), .A2(n575), .B1(data_out[45]), .B2(n569), .ZN(
        n2322) );
  INV_X1 U1029 ( .I(n2320), .ZN(n661) );
  AOI22_X1 U1030 ( .A1(N229), .A2(n575), .B1(data_out[47]), .B2(n569), .ZN(
        n2320) );
  INV_X1 U1031 ( .I(n2325), .ZN(n666) );
  AOI22_X1 U1032 ( .A1(N224), .A2(n575), .B1(data_out[42]), .B2(n569), .ZN(
        n2325) );
  INV_X1 U1033 ( .I(n2331), .ZN(n672) );
  AOI22_X1 U1034 ( .A1(N218), .A2(n575), .B1(data_out[36]), .B2(n569), .ZN(
        n2331) );
  INV_X1 U1035 ( .I(n2329), .ZN(n670) );
  AOI22_X1 U1036 ( .A1(N220), .A2(n575), .B1(data_out[38]), .B2(n569), .ZN(
        n2329) );
  INV_X1 U1037 ( .I(n2323), .ZN(n664) );
  AOI22_X1 U1038 ( .A1(N226), .A2(n575), .B1(data_out[44]), .B2(n569), .ZN(
        n2323) );
  INV_X1 U1039 ( .I(n2321), .ZN(n662) );
  AOI22_X1 U1040 ( .A1(N228), .A2(n575), .B1(data_out[46]), .B2(n569), .ZN(
        n2321) );
  INV_X1 U1041 ( .I(n2319), .ZN(n660) );
  AOI22_X1 U1042 ( .A1(N230), .A2(n576), .B1(data_out[48]), .B2(n570), .ZN(
        n2319) );
  INV_X1 U1043 ( .I(n2318), .ZN(n659) );
  AOI22_X1 U1044 ( .A1(N231), .A2(n576), .B1(data_out[49]), .B2(n570), .ZN(
        n2318) );
  INV_X1 U1045 ( .I(n2317), .ZN(n658) );
  AOI22_X1 U1046 ( .A1(N232), .A2(n576), .B1(data_out[50]), .B2(n570), .ZN(
        n2317) );
  INV_X1 U1047 ( .I(n2316), .ZN(n657) );
  AOI22_X1 U1048 ( .A1(N233), .A2(n576), .B1(data_out[51]), .B2(n570), .ZN(
        n2316) );
  INV_X1 U1049 ( .I(n2315), .ZN(n656) );
  AOI22_X1 U1050 ( .A1(N234), .A2(n576), .B1(data_out[52]), .B2(n570), .ZN(
        n2315) );
  INV_X1 U1051 ( .I(n2314), .ZN(n655) );
  AOI22_X1 U1052 ( .A1(N235), .A2(n576), .B1(data_out[53]), .B2(n570), .ZN(
        n2314) );
  INV_X1 U1053 ( .I(n2313), .ZN(n654) );
  AOI22_X1 U1054 ( .A1(N236), .A2(n576), .B1(data_out[54]), .B2(n570), .ZN(
        n2313) );
  INV_X1 U1055 ( .I(n2312), .ZN(n653) );
  AOI22_X1 U1056 ( .A1(N237), .A2(n576), .B1(data_out[55]), .B2(n570), .ZN(
        n2312) );
  INV_X1 U1057 ( .I(n2311), .ZN(n652) );
  AOI22_X1 U1058 ( .A1(N238), .A2(n576), .B1(data_out[56]), .B2(n570), .ZN(
        n2311) );
  INV_X1 U1059 ( .I(n2310), .ZN(n651) );
  AOI22_X1 U1060 ( .A1(N239), .A2(n576), .B1(data_out[57]), .B2(n570), .ZN(
        n2310) );
  INV_X1 U1061 ( .I(n2309), .ZN(n650) );
  AOI22_X1 U1062 ( .A1(N240), .A2(n576), .B1(data_out[58]), .B2(n570), .ZN(
        n2309) );
  INV_X1 U1063 ( .I(n2308), .ZN(n649) );
  AOI22_X1 U1064 ( .A1(N241), .A2(n576), .B1(data_out[59]), .B2(n570), .ZN(
        n2308) );
  OAI21_X1 U1065 ( .A1(n774), .A2(n478), .B(n2010), .ZN(n1803) );
  NAND2_X1 U1066 ( .A1(rd_ptr[0]), .A2(n2009), .ZN(n2010) );
  INV_X1 U1067 ( .I(n2128), .ZN(n644) );
  AOI22_X1 U1068 ( .A1(n487), .A2(wr_ptr[63]), .B1(n471), .B2(nxt_wr_ptr[63]), 
        .ZN(n2128) );
  INV_X1 U1069 ( .I(n2124), .ZN(n901) );
  AOI22_X1 U1070 ( .A1(n489), .A2(wr_ptr[60]), .B1(n471), .B2(nxt_wr_ptr[60]), 
        .ZN(n2124) );
  INV_X1 U1071 ( .I(n2125), .ZN(n900) );
  AOI22_X1 U1072 ( .A1(n485), .A2(wr_ptr[61]), .B1(n471), .B2(nxt_wr_ptr[61]), 
        .ZN(n2125) );
  INV_X1 U1073 ( .I(n2126), .ZN(n899) );
  AOI22_X1 U1074 ( .A1(n486), .A2(wr_ptr[62]), .B1(n471), .B2(nxt_wr_ptr[62]), 
        .ZN(n2126) );
  INV_X1 U1075 ( .I(full), .ZN(n1712) );
  INV_X1 U1076 ( .I(n2121), .ZN(n904) );
  AOI22_X1 U1077 ( .A1(n486), .A2(wr_ptr[57]), .B1(n470), .B2(nxt_wr_ptr[57]), 
        .ZN(n2121) );
  INV_X1 U1078 ( .I(n2117), .ZN(n908) );
  AOI22_X1 U1079 ( .A1(n489), .A2(wr_ptr[53]), .B1(n470), .B2(nxt_wr_ptr[53]), 
        .ZN(n2117) );
  INV_X1 U1080 ( .I(n2112), .ZN(n912) );
  AOI22_X1 U1081 ( .A1(n489), .A2(wr_ptr[42]), .B1(n470), .B2(nxt_wr_ptr[42]), 
        .ZN(n2112) );
  INV_X1 U1082 ( .I(n2109), .ZN(n915) );
  AOI22_X1 U1083 ( .A1(n489), .A2(wr_ptr[39]), .B1(n469), .B2(nxt_wr_ptr[39]), 
        .ZN(n2109) );
  INV_X1 U1084 ( .I(n2105), .ZN(n919) );
  AOI22_X1 U1085 ( .A1(n489), .A2(wr_ptr[35]), .B1(n469), .B2(nxt_wr_ptr[35]), 
        .ZN(n2105) );
  INV_X1 U1086 ( .I(n2101), .ZN(n923) );
  AOI22_X1 U1087 ( .A1(n488), .A2(wr_ptr[31]), .B1(n469), .B2(nxt_wr_ptr[31]), 
        .ZN(n2101) );
  INV_X1 U1088 ( .I(n2098), .ZN(n926) );
  AOI22_X1 U1089 ( .A1(n488), .A2(wr_ptr[28]), .B1(n468), .B2(nxt_wr_ptr[28]), 
        .ZN(n2098) );
  INV_X1 U1090 ( .I(n2094), .ZN(n930) );
  AOI22_X1 U1091 ( .A1(n488), .A2(wr_ptr[24]), .B1(n468), .B2(nxt_wr_ptr[24]), 
        .ZN(n2094) );
  INV_X1 U1092 ( .I(n2090), .ZN(n934) );
  AOI22_X1 U1093 ( .A1(n488), .A2(wr_ptr[20]), .B1(n468), .B2(nxt_wr_ptr[20]), 
        .ZN(n2090) );
  INV_X1 U1094 ( .I(n2087), .ZN(n937) );
  AOI22_X1 U1095 ( .A1(n488), .A2(wr_ptr[17]), .B1(n468), .B2(nxt_wr_ptr[17]), 
        .ZN(n2087) );
  INV_X1 U1096 ( .I(n2083), .ZN(n941) );
  AOI22_X1 U1097 ( .A1(n487), .A2(wr_ptr[13]), .B1(n467), .B2(nxt_wr_ptr[13]), 
        .ZN(n2083) );
  INV_X1 U1098 ( .I(n2079), .ZN(n945) );
  AOI22_X1 U1099 ( .A1(n487), .A2(wr_ptr[6]), .B1(n467), .B2(nxt_wr_ptr[6]), 
        .ZN(n2079) );
  INV_X1 U1100 ( .I(n2122), .ZN(n903) );
  AOI22_X1 U1101 ( .A1(n489), .A2(wr_ptr[58]), .B1(n470), .B2(nxt_wr_ptr[58]), 
        .ZN(n2122) );
  INV_X1 U1102 ( .I(n2118), .ZN(n907) );
  AOI22_X1 U1103 ( .A1(n489), .A2(wr_ptr[54]), .B1(n470), .B2(nxt_wr_ptr[54]), 
        .ZN(n2118) );
  INV_X1 U1104 ( .I(n2113), .ZN(n911) );
  AOI22_X1 U1105 ( .A1(n489), .A2(wr_ptr[43]), .B1(n470), .B2(nxt_wr_ptr[43]), 
        .ZN(n2113) );
  INV_X1 U1106 ( .I(n2106), .ZN(n918) );
  AOI22_X1 U1107 ( .A1(n489), .A2(wr_ptr[36]), .B1(n469), .B2(nxt_wr_ptr[36]), 
        .ZN(n2106) );
  INV_X1 U1108 ( .I(n2102), .ZN(n922) );
  AOI22_X1 U1109 ( .A1(n489), .A2(wr_ptr[32]), .B1(n469), .B2(nxt_wr_ptr[32]), 
        .ZN(n2102) );
  INV_X1 U1110 ( .I(n2099), .ZN(n925) );
  AOI22_X1 U1111 ( .A1(n488), .A2(wr_ptr[29]), .B1(n469), .B2(nxt_wr_ptr[29]), 
        .ZN(n2099) );
  INV_X1 U1112 ( .I(n2095), .ZN(n929) );
  AOI22_X1 U1113 ( .A1(n488), .A2(wr_ptr[25]), .B1(n468), .B2(nxt_wr_ptr[25]), 
        .ZN(n2095) );
  INV_X1 U1114 ( .I(n2091), .ZN(n933) );
  AOI22_X1 U1115 ( .A1(n488), .A2(wr_ptr[21]), .B1(n468), .B2(nxt_wr_ptr[21]), 
        .ZN(n2091) );
  INV_X1 U1116 ( .I(n2088), .ZN(n936) );
  AOI22_X1 U1117 ( .A1(n488), .A2(wr_ptr[18]), .B1(n468), .B2(nxt_wr_ptr[18]), 
        .ZN(n2088) );
  INV_X1 U1118 ( .I(n2084), .ZN(n940) );
  AOI22_X1 U1119 ( .A1(n487), .A2(wr_ptr[14]), .B1(n467), .B2(nxt_wr_ptr[14]), 
        .ZN(n2084) );
  INV_X1 U1120 ( .I(n2080), .ZN(n944) );
  AOI22_X1 U1121 ( .A1(n487), .A2(wr_ptr[7]), .B1(n467), .B2(nxt_wr_ptr[7]), 
        .ZN(n2080) );
  INV_X1 U1122 ( .I(n2077), .ZN(n947) );
  AOI22_X1 U1123 ( .A1(n487), .A2(wr_ptr[3]), .B1(n467), .B2(nxt_wr_ptr[3]), 
        .ZN(n2077) );
  INV_X1 U1124 ( .I(n2123), .ZN(n902) );
  AOI22_X1 U1125 ( .A1(n488), .A2(wr_ptr[59]), .B1(n470), .B2(nxt_wr_ptr[59]), 
        .ZN(n2123) );
  INV_X1 U1126 ( .I(n2119), .ZN(n906) );
  AOI22_X1 U1127 ( .A1(n485), .A2(wr_ptr[55]), .B1(n470), .B2(nxt_wr_ptr[55]), 
        .ZN(n2119) );
  INV_X1 U1128 ( .I(n2114), .ZN(n910) );
  AOI22_X1 U1129 ( .A1(n489), .A2(wr_ptr[44]), .B1(n470), .B2(nxt_wr_ptr[44]), 
        .ZN(n2114) );
  INV_X1 U1130 ( .I(n2110), .ZN(n914) );
  AOI22_X1 U1131 ( .A1(n489), .A2(wr_ptr[40]), .B1(n469), .B2(nxt_wr_ptr[40]), 
        .ZN(n2110) );
  INV_X1 U1132 ( .I(n2107), .ZN(n917) );
  AOI22_X1 U1133 ( .A1(n489), .A2(wr_ptr[37]), .B1(n469), .B2(nxt_wr_ptr[37]), 
        .ZN(n2107) );
  INV_X1 U1134 ( .I(n2103), .ZN(n921) );
  AOI22_X1 U1135 ( .A1(n489), .A2(wr_ptr[33]), .B1(n469), .B2(nxt_wr_ptr[33]), 
        .ZN(n2103) );
  INV_X1 U1136 ( .I(n2096), .ZN(n928) );
  AOI22_X1 U1137 ( .A1(n488), .A2(wr_ptr[26]), .B1(n468), .B2(nxt_wr_ptr[26]), 
        .ZN(n2096) );
  INV_X1 U1138 ( .I(n2092), .ZN(n932) );
  AOI22_X1 U1139 ( .A1(n488), .A2(wr_ptr[22]), .B1(n468), .B2(nxt_wr_ptr[22]), 
        .ZN(n2092) );
  INV_X1 U1140 ( .I(n2089), .ZN(n935) );
  AOI22_X1 U1141 ( .A1(n488), .A2(wr_ptr[19]), .B1(n468), .B2(nxt_wr_ptr[19]), 
        .ZN(n2089) );
  INV_X1 U1142 ( .I(n2085), .ZN(n939) );
  AOI22_X1 U1143 ( .A1(n488), .A2(wr_ptr[15]), .B1(n467), .B2(nxt_wr_ptr[15]), 
        .ZN(n2085) );
  INV_X1 U1144 ( .I(n2081), .ZN(n943) );
  AOI22_X1 U1145 ( .A1(n487), .A2(wr_ptr[8]), .B1(n467), .B2(nxt_wr_ptr[8]), 
        .ZN(n2081) );
  INV_X1 U1146 ( .I(n2076), .ZN(n948) );
  AOI22_X1 U1147 ( .A1(n487), .A2(wr_ptr[2]), .B1(n467), .B2(nxt_wr_ptr[2]), 
        .ZN(n2076) );
  INV_X1 U1148 ( .I(n2075), .ZN(n949) );
  AOI22_X1 U1149 ( .A1(n487), .A2(wr_ptr[1]), .B1(n467), .B2(nxt_wr_ptr[1]), 
        .ZN(n2075) );
  INV_X1 U1150 ( .I(n2120), .ZN(n905) );
  AOI22_X1 U1151 ( .A1(n485), .A2(wr_ptr[56]), .B1(n470), .B2(nxt_wr_ptr[56]), 
        .ZN(n2120) );
  INV_X1 U1152 ( .I(n2115), .ZN(n909) );
  AOI22_X1 U1153 ( .A1(n489), .A2(wr_ptr[45]), .B1(n470), .B2(nxt_wr_ptr[45]), 
        .ZN(n2115) );
  INV_X1 U1154 ( .I(n2111), .ZN(n913) );
  AOI22_X1 U1155 ( .A1(n489), .A2(wr_ptr[41]), .B1(n470), .B2(nxt_wr_ptr[41]), 
        .ZN(n2111) );
  INV_X1 U1156 ( .I(n2108), .ZN(n916) );
  AOI22_X1 U1157 ( .A1(n489), .A2(wr_ptr[38]), .B1(n469), .B2(nxt_wr_ptr[38]), 
        .ZN(n2108) );
  INV_X1 U1158 ( .I(n2104), .ZN(n920) );
  AOI22_X1 U1159 ( .A1(n489), .A2(wr_ptr[34]), .B1(n469), .B2(nxt_wr_ptr[34]), 
        .ZN(n2104) );
  INV_X1 U1160 ( .I(n2100), .ZN(n924) );
  AOI22_X1 U1161 ( .A1(n488), .A2(wr_ptr[30]), .B1(n469), .B2(nxt_wr_ptr[30]), 
        .ZN(n2100) );
  INV_X1 U1162 ( .I(n2097), .ZN(n927) );
  AOI22_X1 U1163 ( .A1(n488), .A2(wr_ptr[27]), .B1(n468), .B2(nxt_wr_ptr[27]), 
        .ZN(n2097) );
  INV_X1 U1164 ( .I(n2093), .ZN(n931) );
  AOI22_X1 U1165 ( .A1(n488), .A2(wr_ptr[23]), .B1(n468), .B2(nxt_wr_ptr[23]), 
        .ZN(n2093) );
  INV_X1 U1166 ( .I(n2086), .ZN(n938) );
  AOI22_X1 U1167 ( .A1(n488), .A2(wr_ptr[16]), .B1(n467), .B2(nxt_wr_ptr[16]), 
        .ZN(n2086) );
  INV_X1 U1168 ( .I(n2082), .ZN(n942) );
  AOI22_X1 U1169 ( .A1(n487), .A2(wr_ptr[9]), .B1(n467), .B2(nxt_wr_ptr[9]), 
        .ZN(n2082) );
  INV_X1 U1170 ( .I(n2078), .ZN(n946) );
  AOI22_X1 U1171 ( .A1(n487), .A2(wr_ptr[5]), .B1(n467), .B2(nxt_wr_ptr[5]), 
        .ZN(n2078) );
  NAND4_X1 U1172 ( .A1(n2217), .A2(n2216), .A3(wr_ptr[0]), .A4(n2215), .ZN(
        n2281) );
  NOR3_X1 U1173 ( .A1(rst), .A2(wr_ptr[2]), .A3(wr_ptr[1]), .ZN(n2215) );
  INV_X1 U1174 ( .I(n2218), .ZN(n1711) );
  AOI22_X1 U1175 ( .A1(n563), .A2(data_in[0]), .B1(n532), .B2(queue[64]), .ZN(
        n2218) );
  INV_X1 U1176 ( .I(n2219), .ZN(n1710) );
  AOI22_X1 U1177 ( .A1(n563), .A2(data_in[1]), .B1(n532), .B2(queue[65]), .ZN(
        n2219) );
  INV_X1 U1178 ( .I(n2220), .ZN(n1709) );
  AOI22_X1 U1179 ( .A1(n563), .A2(data_in[2]), .B1(n532), .B2(queue[66]), .ZN(
        n2220) );
  INV_X1 U1180 ( .I(n2221), .ZN(n1708) );
  AOI22_X1 U1181 ( .A1(n563), .A2(data_in[3]), .B1(n532), .B2(queue[67]), .ZN(
        n2221) );
  INV_X1 U1182 ( .I(n2222), .ZN(n1707) );
  AOI22_X1 U1183 ( .A1(n562), .A2(data_in[4]), .B1(n532), .B2(queue[68]), .ZN(
        n2222) );
  INV_X1 U1184 ( .I(n2223), .ZN(n1706) );
  AOI22_X1 U1185 ( .A1(n562), .A2(data_in[5]), .B1(n532), .B2(queue[69]), .ZN(
        n2223) );
  INV_X1 U1186 ( .I(n2224), .ZN(n1705) );
  AOI22_X1 U1187 ( .A1(n561), .A2(data_in[6]), .B1(n532), .B2(queue[70]), .ZN(
        n2224) );
  INV_X1 U1188 ( .I(n2225), .ZN(n1704) );
  AOI22_X1 U1189 ( .A1(n561), .A2(data_in[7]), .B1(n532), .B2(queue[71]), .ZN(
        n2225) );
  INV_X1 U1190 ( .I(n2226), .ZN(n1703) );
  AOI22_X1 U1191 ( .A1(n560), .A2(data_in[8]), .B1(n532), .B2(queue[72]), .ZN(
        n2226) );
  INV_X1 U1192 ( .I(n2227), .ZN(n1702) );
  AOI22_X1 U1193 ( .A1(n560), .A2(data_in[9]), .B1(n532), .B2(queue[73]), .ZN(
        n2227) );
  INV_X1 U1194 ( .I(n2228), .ZN(n1701) );
  AOI22_X1 U1195 ( .A1(n559), .A2(data_in[10]), .B1(n532), .B2(queue[74]), 
        .ZN(n2228) );
  INV_X1 U1196 ( .I(n2229), .ZN(n1700) );
  AOI22_X1 U1197 ( .A1(n559), .A2(data_in[11]), .B1(n532), .B2(queue[75]), 
        .ZN(n2229) );
  INV_X1 U1198 ( .I(n2230), .ZN(n1699) );
  AOI22_X1 U1199 ( .A1(n558), .A2(data_in[12]), .B1(n533), .B2(queue[76]), 
        .ZN(n2230) );
  INV_X1 U1200 ( .I(n2231), .ZN(n1698) );
  AOI22_X1 U1201 ( .A1(n558), .A2(data_in[13]), .B1(n533), .B2(queue[77]), 
        .ZN(n2231) );
  INV_X1 U1202 ( .I(n2232), .ZN(n1697) );
  AOI22_X1 U1203 ( .A1(n557), .A2(data_in[14]), .B1(n533), .B2(queue[78]), 
        .ZN(n2232) );
  INV_X1 U1204 ( .I(n2233), .ZN(n1696) );
  AOI22_X1 U1205 ( .A1(n557), .A2(data_in[15]), .B1(n533), .B2(queue[79]), 
        .ZN(n2233) );
  INV_X1 U1206 ( .I(n2234), .ZN(n1695) );
  AOI22_X1 U1207 ( .A1(n556), .A2(data_in[16]), .B1(n533), .B2(queue[80]), 
        .ZN(n2234) );
  INV_X1 U1208 ( .I(n2235), .ZN(n1694) );
  AOI22_X1 U1209 ( .A1(n556), .A2(data_in[17]), .B1(n533), .B2(queue[81]), 
        .ZN(n2235) );
  INV_X1 U1210 ( .I(n2236), .ZN(n1693) );
  AOI22_X1 U1211 ( .A1(n555), .A2(data_in[18]), .B1(n533), .B2(queue[82]), 
        .ZN(n2236) );
  INV_X1 U1212 ( .I(n2237), .ZN(n1692) );
  AOI22_X1 U1213 ( .A1(n555), .A2(data_in[19]), .B1(n533), .B2(queue[83]), 
        .ZN(n2237) );
  INV_X1 U1214 ( .I(n2238), .ZN(n1691) );
  AOI22_X1 U1215 ( .A1(n554), .A2(data_in[20]), .B1(n533), .B2(queue[84]), 
        .ZN(n2238) );
  INV_X1 U1216 ( .I(n2239), .ZN(n1690) );
  AOI22_X1 U1217 ( .A1(n554), .A2(data_in[21]), .B1(n533), .B2(queue[85]), 
        .ZN(n2239) );
  INV_X1 U1218 ( .I(n2240), .ZN(n1689) );
  AOI22_X1 U1219 ( .A1(n553), .A2(data_in[22]), .B1(n533), .B2(queue[86]), 
        .ZN(n2240) );
  INV_X1 U1220 ( .I(n2241), .ZN(n1688) );
  AOI22_X1 U1221 ( .A1(n553), .A2(data_in[23]), .B1(n533), .B2(queue[87]), 
        .ZN(n2241) );
  INV_X1 U1222 ( .I(n2242), .ZN(n1687) );
  AOI22_X1 U1223 ( .A1(n552), .A2(data_in[24]), .B1(n534), .B2(queue[88]), 
        .ZN(n2242) );
  INV_X1 U1224 ( .I(n2243), .ZN(n1686) );
  AOI22_X1 U1225 ( .A1(n552), .A2(data_in[25]), .B1(n534), .B2(queue[89]), 
        .ZN(n2243) );
  INV_X1 U1226 ( .I(n2244), .ZN(n1685) );
  AOI22_X1 U1227 ( .A1(n551), .A2(data_in[26]), .B1(n534), .B2(queue[90]), 
        .ZN(n2244) );
  INV_X1 U1228 ( .I(n2245), .ZN(n1684) );
  AOI22_X1 U1229 ( .A1(n551), .A2(data_in[27]), .B1(n534), .B2(queue[91]), 
        .ZN(n2245) );
  INV_X1 U1230 ( .I(n2246), .ZN(n1683) );
  AOI22_X1 U1231 ( .A1(n550), .A2(data_in[28]), .B1(n534), .B2(queue[92]), 
        .ZN(n2246) );
  INV_X1 U1232 ( .I(n2247), .ZN(n1682) );
  AOI22_X1 U1233 ( .A1(n550), .A2(data_in[29]), .B1(n534), .B2(queue[93]), 
        .ZN(n2247) );
  INV_X1 U1234 ( .I(n2248), .ZN(n1681) );
  AOI22_X1 U1235 ( .A1(n549), .A2(data_in[30]), .B1(n534), .B2(queue[94]), 
        .ZN(n2248) );
  INV_X1 U1236 ( .I(n2249), .ZN(n1680) );
  AOI22_X1 U1237 ( .A1(n549), .A2(data_in[31]), .B1(n534), .B2(queue[95]), 
        .ZN(n2249) );
  INV_X1 U1238 ( .I(n2250), .ZN(n1679) );
  AOI22_X1 U1239 ( .A1(n548), .A2(data_in[32]), .B1(n534), .B2(queue[96]), 
        .ZN(n2250) );
  INV_X1 U1240 ( .I(n2251), .ZN(n1678) );
  AOI22_X1 U1241 ( .A1(n548), .A2(data_in[33]), .B1(n534), .B2(queue[97]), 
        .ZN(n2251) );
  INV_X1 U1242 ( .I(n2252), .ZN(n1677) );
  AOI22_X1 U1243 ( .A1(n547), .A2(data_in[34]), .B1(n534), .B2(queue[98]), 
        .ZN(n2252) );
  INV_X1 U1244 ( .I(n2253), .ZN(n1676) );
  AOI22_X1 U1245 ( .A1(n547), .A2(data_in[35]), .B1(n534), .B2(queue[99]), 
        .ZN(n2253) );
  NAND4_X1 U1246 ( .A1(n2216), .A2(n1736), .A3(n2217), .A4(n2149), .ZN(n2213)
         );
  NOR3_X1 U1247 ( .A1(wr_ptr[0]), .A2(wr_ptr[2]), .A3(wr_ptr[1]), .ZN(n2149)
         );
  INV_X1 U1248 ( .I(n2278), .ZN(n1651) );
  AOI22_X1 U1249 ( .A1(n538), .A2(data_in[60]), .B1(n537), .B2(queue[124]), 
        .ZN(n2278) );
  INV_X1 U1250 ( .I(n2279), .ZN(n1650) );
  AOI22_X1 U1251 ( .A1(n538), .A2(data_in[61]), .B1(n537), .B2(queue[125]), 
        .ZN(n2279) );
  INV_X1 U1252 ( .I(n2280), .ZN(n1649) );
  AOI22_X1 U1253 ( .A1(n538), .A2(data_in[62]), .B1(n537), .B2(queue[126]), 
        .ZN(n2280) );
  INV_X1 U1254 ( .I(n2282), .ZN(n1648) );
  AOI22_X1 U1255 ( .A1(n540), .A2(data_in[63]), .B1(n537), .B2(queue[127]), 
        .ZN(n2282) );
  INV_X1 U1256 ( .I(n2162), .ZN(n1635) );
  AOI22_X1 U1257 ( .A1(data_in[12]), .A2(n524), .B1(n511), .B2(queue[12]), 
        .ZN(n2162) );
  INV_X1 U1258 ( .I(n2163), .ZN(n1634) );
  AOI22_X1 U1259 ( .A1(data_in[13]), .A2(n524), .B1(n510), .B2(queue[13]), 
        .ZN(n2163) );
  INV_X1 U1260 ( .I(n2164), .ZN(n1633) );
  AOI22_X1 U1261 ( .A1(data_in[14]), .A2(n524), .B1(n510), .B2(queue[14]), 
        .ZN(n2164) );
  INV_X1 U1262 ( .I(n2165), .ZN(n1632) );
  AOI22_X1 U1263 ( .A1(data_in[15]), .A2(n524), .B1(n510), .B2(queue[15]), 
        .ZN(n2165) );
  INV_X1 U1264 ( .I(n2166), .ZN(n1631) );
  AOI22_X1 U1265 ( .A1(data_in[16]), .A2(n524), .B1(n509), .B2(queue[16]), 
        .ZN(n2166) );
  INV_X1 U1266 ( .I(n2167), .ZN(n1630) );
  AOI22_X1 U1267 ( .A1(data_in[17]), .A2(n524), .B1(n509), .B2(queue[17]), 
        .ZN(n2167) );
  INV_X1 U1268 ( .I(n2168), .ZN(n1629) );
  AOI22_X1 U1269 ( .A1(data_in[18]), .A2(n524), .B1(n509), .B2(queue[18]), 
        .ZN(n2168) );
  INV_X1 U1270 ( .I(n2169), .ZN(n1628) );
  AOI22_X1 U1271 ( .A1(data_in[19]), .A2(n524), .B1(n508), .B2(queue[19]), 
        .ZN(n2169) );
  INV_X1 U1272 ( .I(n2170), .ZN(n1627) );
  AOI22_X1 U1273 ( .A1(data_in[20]), .A2(n524), .B1(n508), .B2(queue[20]), 
        .ZN(n2170) );
  INV_X1 U1274 ( .I(n2171), .ZN(n1626) );
  AOI22_X1 U1275 ( .A1(data_in[21]), .A2(n524), .B1(n508), .B2(queue[21]), 
        .ZN(n2171) );
  INV_X1 U1276 ( .I(n2172), .ZN(n1625) );
  AOI22_X1 U1277 ( .A1(data_in[22]), .A2(n524), .B1(n507), .B2(queue[22]), 
        .ZN(n2172) );
  INV_X1 U1278 ( .I(n2173), .ZN(n1624) );
  AOI22_X1 U1279 ( .A1(data_in[23]), .A2(n524), .B1(n507), .B2(queue[23]), 
        .ZN(n2173) );
  INV_X1 U1280 ( .I(n2174), .ZN(n1623) );
  AOI22_X1 U1281 ( .A1(data_in[24]), .A2(n524), .B1(n507), .B2(queue[24]), 
        .ZN(n2174) );
  INV_X1 U1282 ( .I(n2175), .ZN(n1622) );
  AOI22_X1 U1283 ( .A1(data_in[25]), .A2(n524), .B1(n506), .B2(queue[25]), 
        .ZN(n2175) );
  INV_X1 U1284 ( .I(n2176), .ZN(n1621) );
  AOI22_X1 U1285 ( .A1(data_in[26]), .A2(n524), .B1(n506), .B2(queue[26]), 
        .ZN(n2176) );
  INV_X1 U1286 ( .I(n2177), .ZN(n1620) );
  AOI22_X1 U1287 ( .A1(data_in[27]), .A2(n524), .B1(n506), .B2(queue[27]), 
        .ZN(n2177) );
  INV_X1 U1288 ( .I(n2178), .ZN(n1619) );
  AOI22_X1 U1289 ( .A1(data_in[28]), .A2(n524), .B1(n505), .B2(queue[28]), 
        .ZN(n2178) );
  INV_X1 U1290 ( .I(n2179), .ZN(n1618) );
  AOI22_X1 U1291 ( .A1(data_in[29]), .A2(n524), .B1(n505), .B2(queue[29]), 
        .ZN(n2179) );
  INV_X1 U1292 ( .I(n2180), .ZN(n1617) );
  AOI22_X1 U1293 ( .A1(data_in[30]), .A2(n524), .B1(n505), .B2(queue[30]), 
        .ZN(n2180) );
  INV_X1 U1294 ( .I(n2181), .ZN(n1616) );
  AOI22_X1 U1295 ( .A1(data_in[31]), .A2(n524), .B1(n504), .B2(queue[31]), 
        .ZN(n2181) );
  INV_X1 U1296 ( .I(n2182), .ZN(n1615) );
  AOI22_X1 U1297 ( .A1(data_in[32]), .A2(n524), .B1(n504), .B2(queue[32]), 
        .ZN(n2182) );
  INV_X1 U1298 ( .I(n2183), .ZN(n1614) );
  AOI22_X1 U1299 ( .A1(data_in[33]), .A2(n524), .B1(n504), .B2(queue[33]), 
        .ZN(n2183) );
  INV_X1 U1300 ( .I(n2184), .ZN(n1613) );
  AOI22_X1 U1301 ( .A1(data_in[34]), .A2(n524), .B1(n503), .B2(queue[34]), 
        .ZN(n2184) );
  INV_X1 U1302 ( .I(n2185), .ZN(n1612) );
  AOI22_X1 U1303 ( .A1(data_in[35]), .A2(n524), .B1(n503), .B2(queue[35]), 
        .ZN(n2185) );
  INV_X1 U1304 ( .I(n2254), .ZN(n1675) );
  AOI22_X1 U1305 ( .A1(n546), .A2(data_in[36]), .B1(n535), .B2(queue[100]), 
        .ZN(n2254) );
  INV_X1 U1306 ( .I(n2255), .ZN(n1674) );
  AOI22_X1 U1307 ( .A1(n546), .A2(data_in[37]), .B1(n535), .B2(queue[101]), 
        .ZN(n2255) );
  INV_X1 U1308 ( .I(n2256), .ZN(n1673) );
  AOI22_X1 U1309 ( .A1(n545), .A2(data_in[38]), .B1(n535), .B2(queue[102]), 
        .ZN(n2256) );
  INV_X1 U1310 ( .I(n2257), .ZN(n1672) );
  AOI22_X1 U1311 ( .A1(n545), .A2(data_in[39]), .B1(n535), .B2(queue[103]), 
        .ZN(n2257) );
  INV_X1 U1312 ( .I(n2258), .ZN(n1671) );
  AOI22_X1 U1313 ( .A1(n544), .A2(data_in[40]), .B1(n535), .B2(queue[104]), 
        .ZN(n2258) );
  INV_X1 U1314 ( .I(n2259), .ZN(n1670) );
  AOI22_X1 U1315 ( .A1(n544), .A2(data_in[41]), .B1(n535), .B2(queue[105]), 
        .ZN(n2259) );
  INV_X1 U1316 ( .I(n2260), .ZN(n1669) );
  AOI22_X1 U1317 ( .A1(n547), .A2(data_in[42]), .B1(n535), .B2(queue[106]), 
        .ZN(n2260) );
  INV_X1 U1318 ( .I(n2261), .ZN(n1668) );
  AOI22_X1 U1319 ( .A1(n546), .A2(data_in[43]), .B1(n535), .B2(queue[107]), 
        .ZN(n2261) );
  INV_X1 U1320 ( .I(n2262), .ZN(n1667) );
  AOI22_X1 U1321 ( .A1(n543), .A2(data_in[44]), .B1(n535), .B2(queue[108]), 
        .ZN(n2262) );
  INV_X1 U1322 ( .I(n2263), .ZN(n1666) );
  AOI22_X1 U1323 ( .A1(n543), .A2(data_in[45]), .B1(n535), .B2(queue[109]), 
        .ZN(n2263) );
  INV_X1 U1324 ( .I(n2264), .ZN(n1665) );
  AOI22_X1 U1325 ( .A1(n542), .A2(data_in[46]), .B1(n535), .B2(queue[110]), 
        .ZN(n2264) );
  INV_X1 U1326 ( .I(n2265), .ZN(n1664) );
  AOI22_X1 U1327 ( .A1(n542), .A2(data_in[47]), .B1(n535), .B2(queue[111]), 
        .ZN(n2265) );
  INV_X1 U1328 ( .I(n2266), .ZN(n1663) );
  AOI22_X1 U1329 ( .A1(n541), .A2(data_in[48]), .B1(n536), .B2(queue[112]), 
        .ZN(n2266) );
  INV_X1 U1330 ( .I(n2267), .ZN(n1662) );
  AOI22_X1 U1331 ( .A1(n541), .A2(data_in[49]), .B1(n536), .B2(queue[113]), 
        .ZN(n2267) );
  INV_X1 U1332 ( .I(n2268), .ZN(n1661) );
  AOI22_X1 U1333 ( .A1(n541), .A2(data_in[50]), .B1(n536), .B2(queue[114]), 
        .ZN(n2268) );
  INV_X1 U1334 ( .I(n2269), .ZN(n1660) );
  AOI22_X1 U1335 ( .A1(n541), .A2(data_in[51]), .B1(n536), .B2(queue[115]), 
        .ZN(n2269) );
  INV_X1 U1336 ( .I(n2270), .ZN(n1659) );
  AOI22_X1 U1337 ( .A1(n543), .A2(data_in[52]), .B1(n536), .B2(queue[116]), 
        .ZN(n2270) );
  INV_X1 U1338 ( .I(n2271), .ZN(n1658) );
  AOI22_X1 U1339 ( .A1(n542), .A2(data_in[53]), .B1(n536), .B2(queue[117]), 
        .ZN(n2271) );
  INV_X1 U1340 ( .I(n2272), .ZN(n1657) );
  AOI22_X1 U1341 ( .A1(n540), .A2(data_in[54]), .B1(n536), .B2(queue[118]), 
        .ZN(n2272) );
  INV_X1 U1342 ( .I(n2273), .ZN(n1656) );
  AOI22_X1 U1343 ( .A1(n540), .A2(data_in[55]), .B1(n536), .B2(queue[119]), 
        .ZN(n2273) );
  INV_X1 U1344 ( .I(n2274), .ZN(n1655) );
  AOI22_X1 U1345 ( .A1(n539), .A2(data_in[56]), .B1(n536), .B2(queue[120]), 
        .ZN(n2274) );
  INV_X1 U1346 ( .I(n2275), .ZN(n1654) );
  AOI22_X1 U1347 ( .A1(n539), .A2(data_in[57]), .B1(n536), .B2(queue[121]), 
        .ZN(n2275) );
  INV_X1 U1348 ( .I(n2276), .ZN(n1653) );
  AOI22_X1 U1349 ( .A1(n539), .A2(data_in[58]), .B1(n536), .B2(queue[122]), 
        .ZN(n2276) );
  INV_X1 U1350 ( .I(n2277), .ZN(n1652) );
  AOI22_X1 U1351 ( .A1(n538), .A2(data_in[59]), .B1(n536), .B2(queue[123]), 
        .ZN(n2277) );
  INV_X1 U1352 ( .I(n2150), .ZN(n1647) );
  AOI22_X1 U1353 ( .A1(data_in[0]), .A2(n524), .B1(n515), .B2(queue[0]), .ZN(
        n2150) );
  INV_X1 U1354 ( .I(n2210), .ZN(n954) );
  AOI22_X1 U1355 ( .A1(data_in[60]), .A2(n524), .B1(n495), .B2(queue[60]), 
        .ZN(n2210) );
  INV_X1 U1356 ( .I(n2211), .ZN(n953) );
  AOI22_X1 U1357 ( .A1(data_in[61]), .A2(n524), .B1(n494), .B2(queue[61]), 
        .ZN(n2211) );
  INV_X1 U1358 ( .I(n2212), .ZN(n952) );
  AOI22_X1 U1359 ( .A1(data_in[62]), .A2(n524), .B1(n494), .B2(queue[62]), 
        .ZN(n2212) );
  INV_X1 U1360 ( .I(n2214), .ZN(n951) );
  AOI22_X1 U1361 ( .A1(data_in[63]), .A2(n524), .B1(n494), .B2(queue[63]), 
        .ZN(n2214) );
  INV_X1 U1362 ( .I(n2151), .ZN(n1646) );
  AOI22_X1 U1363 ( .A1(data_in[1]), .A2(n524), .B1(n514), .B2(queue[1]), .ZN(
        n2151) );
  INV_X1 U1364 ( .I(n2152), .ZN(n1645) );
  AOI22_X1 U1365 ( .A1(data_in[2]), .A2(n524), .B1(n514), .B2(queue[2]), .ZN(
        n2152) );
  INV_X1 U1366 ( .I(n2153), .ZN(n1644) );
  AOI22_X1 U1367 ( .A1(data_in[3]), .A2(n524), .B1(n514), .B2(queue[3]), .ZN(
        n2153) );
  INV_X1 U1368 ( .I(n2154), .ZN(n1643) );
  AOI22_X1 U1369 ( .A1(data_in[4]), .A2(n524), .B1(n513), .B2(queue[4]), .ZN(
        n2154) );
  INV_X1 U1370 ( .I(n2155), .ZN(n1642) );
  AOI22_X1 U1371 ( .A1(data_in[5]), .A2(n524), .B1(n513), .B2(queue[5]), .ZN(
        n2155) );
  INV_X1 U1372 ( .I(n2156), .ZN(n1641) );
  AOI22_X1 U1373 ( .A1(data_in[6]), .A2(n524), .B1(n513), .B2(queue[6]), .ZN(
        n2156) );
  INV_X1 U1374 ( .I(n2157), .ZN(n1640) );
  AOI22_X1 U1375 ( .A1(data_in[7]), .A2(n524), .B1(n512), .B2(queue[7]), .ZN(
        n2157) );
  INV_X1 U1376 ( .I(n2158), .ZN(n1639) );
  AOI22_X1 U1377 ( .A1(data_in[8]), .A2(n524), .B1(n512), .B2(queue[8]), .ZN(
        n2158) );
  INV_X1 U1378 ( .I(n2159), .ZN(n1638) );
  AOI22_X1 U1379 ( .A1(data_in[9]), .A2(n524), .B1(n512), .B2(queue[9]), .ZN(
        n2159) );
  INV_X1 U1380 ( .I(n2160), .ZN(n1637) );
  AOI22_X1 U1381 ( .A1(data_in[10]), .A2(n524), .B1(n511), .B2(queue[10]), 
        .ZN(n2160) );
  INV_X1 U1382 ( .I(n2161), .ZN(n1636) );
  AOI22_X1 U1383 ( .A1(data_in[11]), .A2(n524), .B1(n511), .B2(queue[11]), 
        .ZN(n2161) );
  INV_X1 U1384 ( .I(n2186), .ZN(n1611) );
  AOI22_X1 U1385 ( .A1(data_in[36]), .A2(n524), .B1(n503), .B2(queue[36]), 
        .ZN(n2186) );
  INV_X1 U1386 ( .I(n2187), .ZN(n1336) );
  AOI22_X1 U1387 ( .A1(data_in[37]), .A2(n524), .B1(n502), .B2(queue[37]), 
        .ZN(n2187) );
  INV_X1 U1388 ( .I(n2188), .ZN(n976) );
  AOI22_X1 U1389 ( .A1(data_in[38]), .A2(n524), .B1(n502), .B2(queue[38]), 
        .ZN(n2188) );
  INV_X1 U1390 ( .I(n2189), .ZN(n975) );
  AOI22_X1 U1391 ( .A1(data_in[39]), .A2(n524), .B1(n502), .B2(queue[39]), 
        .ZN(n2189) );
  INV_X1 U1392 ( .I(n2190), .ZN(n974) );
  AOI22_X1 U1393 ( .A1(data_in[40]), .A2(n524), .B1(n501), .B2(queue[40]), 
        .ZN(n2190) );
  INV_X1 U1394 ( .I(n2191), .ZN(n973) );
  AOI22_X1 U1395 ( .A1(data_in[41]), .A2(n524), .B1(n501), .B2(queue[41]), 
        .ZN(n2191) );
  INV_X1 U1396 ( .I(n2192), .ZN(n972) );
  AOI22_X1 U1397 ( .A1(data_in[42]), .A2(n524), .B1(n501), .B2(queue[42]), 
        .ZN(n2192) );
  INV_X1 U1398 ( .I(n2193), .ZN(n971) );
  AOI22_X1 U1399 ( .A1(data_in[43]), .A2(n524), .B1(n500), .B2(queue[43]), 
        .ZN(n2193) );
  INV_X1 U1400 ( .I(n2194), .ZN(n970) );
  AOI22_X1 U1401 ( .A1(data_in[44]), .A2(n524), .B1(n500), .B2(queue[44]), 
        .ZN(n2194) );
  INV_X1 U1402 ( .I(n2195), .ZN(n969) );
  AOI22_X1 U1403 ( .A1(data_in[45]), .A2(n524), .B1(n500), .B2(queue[45]), 
        .ZN(n2195) );
  INV_X1 U1404 ( .I(n2196), .ZN(n968) );
  AOI22_X1 U1405 ( .A1(data_in[46]), .A2(n524), .B1(n499), .B2(queue[46]), 
        .ZN(n2196) );
  INV_X1 U1406 ( .I(n2197), .ZN(n967) );
  AOI22_X1 U1407 ( .A1(data_in[47]), .A2(n524), .B1(n499), .B2(queue[47]), 
        .ZN(n2197) );
  INV_X1 U1408 ( .I(n2198), .ZN(n966) );
  AOI22_X1 U1409 ( .A1(data_in[48]), .A2(n524), .B1(n499), .B2(queue[48]), 
        .ZN(n2198) );
  INV_X1 U1410 ( .I(n2199), .ZN(n965) );
  AOI22_X1 U1411 ( .A1(data_in[49]), .A2(n524), .B1(n498), .B2(queue[49]), 
        .ZN(n2199) );
  INV_X1 U1412 ( .I(n2200), .ZN(n964) );
  AOI22_X1 U1413 ( .A1(data_in[50]), .A2(n524), .B1(n498), .B2(queue[50]), 
        .ZN(n2200) );
  INV_X1 U1414 ( .I(n2201), .ZN(n963) );
  AOI22_X1 U1415 ( .A1(data_in[51]), .A2(n524), .B1(n498), .B2(queue[51]), 
        .ZN(n2201) );
  INV_X1 U1416 ( .I(n2202), .ZN(n962) );
  AOI22_X1 U1417 ( .A1(data_in[52]), .A2(n524), .B1(n497), .B2(queue[52]), 
        .ZN(n2202) );
  INV_X1 U1418 ( .I(n2203), .ZN(n961) );
  AOI22_X1 U1419 ( .A1(data_in[53]), .A2(n524), .B1(n497), .B2(queue[53]), 
        .ZN(n2203) );
  INV_X1 U1420 ( .I(n2204), .ZN(n960) );
  AOI22_X1 U1421 ( .A1(data_in[54]), .A2(n524), .B1(n497), .B2(queue[54]), 
        .ZN(n2204) );
  INV_X1 U1422 ( .I(n2205), .ZN(n959) );
  AOI22_X1 U1423 ( .A1(data_in[55]), .A2(n524), .B1(n496), .B2(queue[55]), 
        .ZN(n2205) );
  INV_X1 U1424 ( .I(n2206), .ZN(n958) );
  AOI22_X1 U1425 ( .A1(data_in[56]), .A2(n524), .B1(n496), .B2(queue[56]), 
        .ZN(n2206) );
  INV_X1 U1426 ( .I(n2207), .ZN(n957) );
  AOI22_X1 U1427 ( .A1(data_in[57]), .A2(n524), .B1(n496), .B2(queue[57]), 
        .ZN(n2207) );
  INV_X1 U1428 ( .I(n2208), .ZN(n956) );
  AOI22_X1 U1429 ( .A1(data_in[58]), .A2(n524), .B1(n495), .B2(queue[58]), 
        .ZN(n2208) );
  INV_X1 U1430 ( .I(n2209), .ZN(n955) );
  AOI22_X1 U1431 ( .A1(data_in[59]), .A2(n524), .B1(n495), .B2(queue[59]), 
        .ZN(n2209) );
  INV_X1 U1432 ( .I(empty), .ZN(n710) );
  OAI22_X1 U1433 ( .A1(n491), .A2(n643), .B1(n487), .B2(n1898), .ZN(n1737) );
  AOI21_X1 U1434 ( .A1(N532), .A2(n1899), .B(rst), .ZN(n1898) );
  INV_X1 U1435 ( .I(rd_ptr[56]), .ZN(n885) );
  OAI22_X1 U1436 ( .A1(n774), .A2(n457), .B1(n2009), .B2(n2007), .ZN(n1740) );
  AOI21_X1 U1437 ( .A1(N246), .A2(n2006), .B(rst), .ZN(n2007) );
  NOR4_X1 U1438 ( .A1(n2137), .A2(n2136), .A3(n2135), .A4(n2134), .ZN(n2148)
         );
  NOR4_X1 U1439 ( .A1(n2146), .A2(n2145), .A3(n2144), .A4(n2143), .ZN(n2147)
         );
  INV_X1 U1440 ( .I(rd_ptr[5]), .ZN(n783) );
  INV_X1 U1441 ( .I(rd_ptr[63]), .ZN(n898) );
  INV_X1 U1442 ( .I(rd_ptr[41]), .ZN(n855) );
  INV_X1 U1443 ( .I(rd_ptr[45]), .ZN(n863) );
  INV_X1 U1444 ( .I(rd_ptr[49]), .ZN(n871) );
  INV_X1 U1445 ( .I(rd_ptr[26]), .ZN(n825) );
  INV_X1 U1446 ( .I(rd_ptr[30]), .ZN(n833) );
  INV_X1 U1447 ( .I(rd_ptr[54]), .ZN(n881) );
  INV_X1 U1448 ( .I(rd_ptr[58]), .ZN(n889) );
  INV_X1 U1449 ( .I(rd_ptr[3]), .ZN(n779) );
  INV_X1 U1450 ( .I(rd_ptr[55]), .ZN(n883) );
  INV_X1 U1451 ( .I(rd_ptr[59]), .ZN(n891) );
  INV_X1 U1452 ( .I(rd_ptr[62]), .ZN(n897) );
  INV_X1 U1453 ( .I(rd_ptr[40]), .ZN(n853) );
  INV_X1 U1454 ( .I(rd_ptr[44]), .ZN(n861) );
  INV_X1 U1455 ( .I(rd_ptr[25]), .ZN(n823) );
  OAI22_X1 U1456 ( .A1(n1713), .A2(n490), .B1(n456), .B2(n643), .ZN(n1866) );
  INV_X1 U1457 ( .I(wr_ptr[0]), .ZN(n1713) );
  INV_X1 U1458 ( .I(rd_ptr[53]), .ZN(n879) );
  INV_X1 U1459 ( .I(rd_ptr[57]), .ZN(n887) );
  INV_X1 U1460 ( .I(rd_ptr[39]), .ZN(n851) );
  INV_X1 U1461 ( .I(rd_ptr[42]), .ZN(n857) );
  INV_X1 U1462 ( .I(rd_ptr[9]), .ZN(n791) );
  INV_X1 U1463 ( .I(rd_ptr[52]), .ZN(n877) );
  INV_X1 U1464 ( .I(rd_ptr[34]), .ZN(n841) );
  INV_X1 U1465 ( .I(rd_ptr[38]), .ZN(n849) );
  INV_X1 U1466 ( .I(rd_ptr[14]), .ZN(n801) );
  INV_X1 U1467 ( .I(rd_ptr[18]), .ZN(n809) );
  INV_X1 U1468 ( .I(rd_ptr[61]), .ZN(n895) );
  INV_X1 U1469 ( .I(rd_ptr[43]), .ZN(n859) );
  INV_X1 U1470 ( .I(rd_ptr[47]), .ZN(n867) );
  INV_X1 U1471 ( .I(rd_ptr[24]), .ZN(n821) );
  INV_X1 U1472 ( .I(rd_ptr[28]), .ZN(n829) );
  INV_X1 U1473 ( .I(rd_ptr[32]), .ZN(n837) );
  INV_X1 U1474 ( .I(rd_ptr[8]), .ZN(n789) );
  INV_X1 U1475 ( .I(rd_ptr[48]), .ZN(n869) );
  INV_X1 U1476 ( .I(rd_ptr[51]), .ZN(n875) );
  INV_X1 U1477 ( .I(rd_ptr[29]), .ZN(n831) );
  INV_X1 U1478 ( .I(rd_ptr[33]), .ZN(n839) );
  INV_X1 U1479 ( .I(rd_ptr[13]), .ZN(n799) );
  INV_X1 U1480 ( .I(rd_ptr[17]), .ZN(n807) );
  NAND3_X1 U1481 ( .A1(n710), .A2(n793), .A3(rd), .ZN(n2283) );
  INV_X1 U1482 ( .I(rd_ptr[60]), .ZN(n893) );
  INV_X1 U1483 ( .I(rd_ptr[6]), .ZN(n785) );
  INV_X1 U1484 ( .I(rd_ptr[46]), .ZN(n865) );
  INV_X1 U1485 ( .I(rd_ptr[23]), .ZN(n819) );
  INV_X1 U1486 ( .I(rd_ptr[27]), .ZN(n827) );
  INV_X1 U1487 ( .I(rd_ptr[31]), .ZN(n835) );
  INV_X1 U1488 ( .I(rd_ptr[11]), .ZN(n795) );
  INV_X1 U1489 ( .I(rd_ptr[22]), .ZN(n817) );
  INV_X1 U1490 ( .I(rd_ptr[7]), .ZN(n787) );
  INV_X1 U1491 ( .I(rd_ptr[50]), .ZN(n873) );
  INV_X1 U1492 ( .I(rd_ptr[36]), .ZN(n845) );
  INV_X1 U1493 ( .I(rd_ptr[12]), .ZN(n797) );
  INV_X1 U1494 ( .I(rd_ptr[16]), .ZN(n805) );
  INV_X1 U1495 ( .I(rd_ptr[37]), .ZN(n847) );
  INV_X1 U1496 ( .I(rd_ptr[21]), .ZN(n815) );
  INV_X1 U1497 ( .I(rd_ptr[10]), .ZN(n793) );
  INV_X1 U1498 ( .I(rd_ptr[4]), .ZN(n781) );
  INV_X1 U1499 ( .I(rd_ptr[35]), .ZN(n843) );
  INV_X1 U1500 ( .I(rd_ptr[15]), .ZN(n803) );
  INV_X1 U1501 ( .I(rd_ptr[20]), .ZN(n813) );
  NAND4_X1 U1502 ( .A1(n1719), .A2(n1721), .A3(n1717), .A4(n2133), .ZN(n2136)
         );
  NOR4_X1 U1503 ( .A1(wr_ptr[16]), .A2(wr_ptr[15]), .A3(wr_ptr[14]), .A4(
        wr_ptr[13]), .ZN(n2133) );
  INV_X1 U1504 ( .I(rd_ptr[19]), .ZN(n811) );
  NOR4_X1 U1505 ( .A1(wr_ptr[9]), .A2(wr_ptr[8]), .A3(wr_ptr[7]), .A4(
        wr_ptr[6]), .ZN(n2138) );
  NOR4_X1 U1506 ( .A1(wr_ptr[39]), .A2(wr_ptr[38]), .A3(wr_ptr[37]), .A4(
        wr_ptr[36]), .ZN(n2129) );
  NAND4_X1 U1507 ( .A1(n2141), .A2(n2140), .A3(n2139), .A4(n2138), .ZN(n2146)
         );
  NOR4_X1 U1508 ( .A1(wr_ptr[56]), .A2(wr_ptr[55]), .A3(wr_ptr[54]), .A4(
        wr_ptr[53]), .ZN(n2141) );
  NOR4_X1 U1509 ( .A1(wr_ptr[5]), .A2(wr_ptr[59]), .A3(wr_ptr[58]), .A4(
        wr_ptr[57]), .ZN(n2140) );
  NOR4_X1 U1510 ( .A1(wr_ptr[63]), .A2(wr_ptr[62]), .A3(wr_ptr[61]), .A4(
        wr_ptr[60]), .ZN(n2139) );
  NAND4_X1 U1511 ( .A1(n2132), .A2(n2131), .A3(n2130), .A4(n2129), .ZN(n2137)
         );
  NOR3_X1 U1512 ( .A1(wr_ptr[25]), .A2(wr_ptr[27]), .A3(wr_ptr[26]), .ZN(n2132) );
  NOR4_X1 U1513 ( .A1(wr_ptr[31]), .A2(wr_ptr[30]), .A3(wr_ptr[29]), .A4(
        wr_ptr[28]), .ZN(n2131) );
  NOR4_X1 U1514 ( .A1(wr_ptr[35]), .A2(wr_ptr[34]), .A3(wr_ptr[33]), .A4(
        wr_ptr[32]), .ZN(n2130) );
  INV_X1 U1515 ( .I(wr_ptr[49]), .ZN(n1729) );
  INV_X1 U1516 ( .I(wr_ptr[52]), .ZN(n1735) );
  INV_X1 U1517 ( .I(wr_ptr[47]), .ZN(n1725) );
  INV_X1 U1518 ( .I(wr_ptr[50]), .ZN(n1731) );
  INV_X1 U1519 ( .I(wr_ptr[48]), .ZN(n1727) );
  INV_X1 U1520 ( .I(wr_ptr[51]), .ZN(n1733) );
  INV_X1 U1521 ( .I(wr_ptr[10]), .ZN(n1717) );
  INV_X1 U1522 ( .I(wr_ptr[46]), .ZN(n1723) );
  INV_X1 U1523 ( .I(wr_ptr[4]), .ZN(n1715) );
  INV_X1 U1524 ( .I(wr_ptr[12]), .ZN(n1721) );
  INV_X1 U1525 ( .I(wr_ptr[11]), .ZN(n1719) );
  NOR4_X1 U1526 ( .A1(n1893), .A2(n1892), .A3(n1891), .A4(n1890), .ZN(n1894)
         );
  NAND4_X1 U1527 ( .A1(nxt_wr_ptr[0]), .A2(n1716), .A3(n1718), .A4(n1720), 
        .ZN(n1878) );
  INV_X1 U1614 ( .I(nxt_wr_ptr[49]), .ZN(n1728) );
  INV_X1 U1615 ( .I(nxt_wr_ptr[12]), .ZN(n1720) );
  INV_X1 U1616 ( .I(nxt_wr_ptr[48]), .ZN(n1726) );
  INV_X1 U1617 ( .I(nxt_wr_ptr[11]), .ZN(n1718) );
  INV_X1 U1618 ( .I(nxt_wr_ptr[46]), .ZN(n1722) );
  INV_X1 U1619 ( .I(nxt_wr_ptr[47]), .ZN(n1724) );
  INV_X1 U1620 ( .I(nxt_wr_ptr[50]), .ZN(n1730) );
  INV_X1 U1621 ( .I(nxt_wr_ptr[10]), .ZN(n1716) );
  INV_X1 U1622 ( .I(nxt_wr_ptr[52]), .ZN(n1734) );
  INV_X1 U1623 ( .I(nxt_wr_ptr[51]), .ZN(n1732) );
  INV_X1 U1624 ( .I(nxt_wr_ptr[4]), .ZN(n1714) );
  INV_X1 U1625 ( .I(nxt_rd_ptr[63]), .ZN(n775) );
  INV_X1 U1626 ( .I(nxt_rd_ptr[5]), .ZN(n782) );
  INV_X1 U1627 ( .I(nxt_rd_ptr[56]), .ZN(n884) );
  INV_X1 U1628 ( .I(nxt_rd_ptr[41]), .ZN(n854) );
  INV_X1 U1629 ( .I(nxt_rd_ptr[55]), .ZN(n882) );
  NAND4_X1 U1630 ( .A1(nxt_rd_ptr[0]), .A2(n792), .A3(n794), .A4(n796), .ZN(
        n1986) );
  INV_X1 U1631 ( .I(nxt_rd_ptr[27]), .ZN(n826) );
  INV_X1 U1632 ( .I(nxt_rd_ptr[12]), .ZN(n796) );
  INV_X1 U1633 ( .I(nxt_rd_ptr[49]), .ZN(n870) );
  INV_X1 U1634 ( .I(nxt_rd_ptr[34]), .ZN(n840) );
  INV_X1 U1635 ( .I(nxt_rd_ptr[45]), .ZN(n862) );
  INV_X1 U1636 ( .I(nxt_rd_ptr[30]), .ZN(n832) );
  INV_X1 U1637 ( .I(nxt_rd_ptr[11]), .ZN(n794) );
  INV_X1 U1638 ( .I(nxt_rd_ptr[48]), .ZN(n868) );
  INV_X1 U1639 ( .I(nxt_rd_ptr[62]), .ZN(n896) );
  INV_X1 U1640 ( .I(nxt_rd_ptr[59]), .ZN(n890) );
  INV_X1 U1641 ( .I(nxt_rd_ptr[33]), .ZN(n838) );
  INV_X1 U1642 ( .I(nxt_rd_ptr[40]), .ZN(n852) );
  INV_X1 U1643 ( .I(nxt_rd_ptr[44]), .ZN(n860) );
  INV_X1 U1644 ( .I(nxt_rd_ptr[26]), .ZN(n824) );
  INV_X1 U1645 ( .I(nxt_rd_ptr[43]), .ZN(n858) );
  INV_X1 U1646 ( .I(nxt_rd_ptr[3]), .ZN(n778) );
  INV_X1 U1647 ( .I(nxt_rd_ptr[54]), .ZN(n880) );
  INV_X1 U1648 ( .I(nxt_rd_ptr[61]), .ZN(n894) );
  INV_X1 U1649 ( .I(nxt_rd_ptr[58]), .ZN(n888) );
  INV_X1 U1650 ( .I(nxt_rd_ptr[25]), .ZN(n822) );
  INV_X1 U1651 ( .I(nxt_rd_ptr[29]), .ZN(n830) );
  INV_X1 U1652 ( .I(nxt_rd_ptr[53]), .ZN(n878) );
  INV_X1 U1653 ( .I(nxt_rd_ptr[9]), .ZN(n790) );
  INV_X1 U1654 ( .I(nxt_rd_ptr[52]), .ZN(n876) );
  INV_X1 U1655 ( .I(nxt_rd_ptr[38]), .ZN(n848) );
  INV_X1 U1656 ( .I(nxt_rd_ptr[16]), .ZN(n804) );
  INV_X1 U1657 ( .I(nxt_rd_ptr[51]), .ZN(n874) );
  INV_X1 U1658 ( .I(nxt_rd_ptr[15]), .ZN(n802) );
  INV_X1 U1659 ( .I(nxt_rd_ptr[19]), .ZN(n810) );
  INV_X1 U1660 ( .I(nxt_rd_ptr[8]), .ZN(n788) );
  INV_X1 U1661 ( .I(nxt_rd_ptr[37]), .ZN(n846) );
  INV_X1 U1662 ( .I(nxt_rd_ptr[47]), .ZN(n866) );
  INV_X1 U1663 ( .I(nxt_rd_ptr[10]), .ZN(n792) );
  INV_X1 U1664 ( .I(nxt_rd_ptr[14]), .ZN(n800) );
  INV_X1 U1665 ( .I(nxt_rd_ptr[7]), .ZN(n786) );
  INV_X1 U1666 ( .I(nxt_rd_ptr[50]), .ZN(n872) );
  INV_X1 U1667 ( .I(nxt_rd_ptr[32]), .ZN(n836) );
  INV_X1 U1668 ( .I(nxt_rd_ptr[18]), .ZN(n808) );
  INV_X1 U1669 ( .I(nxt_rd_ptr[39]), .ZN(n850) );
  INV_X1 U1670 ( .I(nxt_rd_ptr[31]), .ZN(n834) );
  INV_X1 U1671 ( .I(nxt_rd_ptr[60]), .ZN(n892) );
  INV_X1 U1672 ( .I(nxt_rd_ptr[57]), .ZN(n886) );
  INV_X1 U1673 ( .I(nxt_rd_ptr[42]), .ZN(n856) );
  INV_X1 U1674 ( .I(nxt_rd_ptr[46]), .ZN(n864) );
  INV_X1 U1675 ( .I(nxt_rd_ptr[24]), .ZN(n820) );
  INV_X1 U1676 ( .I(nxt_rd_ptr[28]), .ZN(n828) );
  INV_X1 U1677 ( .I(nxt_rd_ptr[2]), .ZN(n777) );
  INV_X1 U1678 ( .I(nxt_rd_ptr[23]), .ZN(n818) );
  INV_X1 U1679 ( .I(nxt_rd_ptr[22]), .ZN(n816) );
  INV_X1 U1680 ( .I(nxt_rd_ptr[36]), .ZN(n844) );
  INV_X1 U1681 ( .I(nxt_rd_ptr[21]), .ZN(n814) );
  INV_X1 U1682 ( .I(nxt_rd_ptr[4]), .ZN(n780) );
  INV_X1 U1683 ( .I(nxt_rd_ptr[35]), .ZN(n842) );
  INV_X1 U1684 ( .I(nxt_rd_ptr[13]), .ZN(n798) );
  INV_X1 U1685 ( .I(nxt_rd_ptr[6]), .ZN(n784) );
  INV_X1 U1686 ( .I(nxt_rd_ptr[17]), .ZN(n806) );
  INV_X1 U1687 ( .I(nxt_rd_ptr[1]), .ZN(n776) );
  INV_X1 U1688 ( .I(nxt_rd_ptr[20]), .ZN(n812) );
  NAND4_X1 U1689 ( .A1(n1916), .A2(n1915), .A3(n1914), .A4(n1913), .ZN(n1917)
         );
  INV_X1 U1690 ( .I(nxt_rd_ptr[0]), .ZN(n774) );
  NAND4_X1 U1691 ( .A1(n1936), .A2(n1935), .A3(n1934), .A4(n1933), .ZN(n1937)
         );
  NAND4_X1 U1692 ( .A1(n1956), .A2(n1955), .A3(n1954), .A4(n1953), .ZN(n1957)
         );
  NAND4_X1 U1693 ( .A1(n1976), .A2(n1975), .A3(n1974), .A4(n1973), .ZN(n1977)
         );
  NAND4_X1 U1694 ( .A1(n1952), .A2(n1951), .A3(n1950), .A4(n1949), .ZN(n1958)
         );
  NAND4_X1 U1695 ( .A1(n1972), .A2(n1971), .A3(n1970), .A4(n1969), .ZN(n1978)
         );
  NAND4_X1 U1696 ( .A1(n1964), .A2(n1963), .A3(n1962), .A4(n1961), .ZN(n1980)
         );
  NAND4_X1 U1697 ( .A1(n1932), .A2(n1931), .A3(n1930), .A4(n1929), .ZN(n1938)
         );
  NAND4_X1 U1698 ( .A1(n1968), .A2(n1967), .A3(n1966), .A4(n1965), .ZN(n1979)
         );
  NAND4_X1 U1699 ( .A1(n1948), .A2(n1947), .A3(n1946), .A4(n1945), .ZN(n1959)
         );
  NAND4_X1 U1700 ( .A1(n1928), .A2(n1927), .A3(n1926), .A4(n1925), .ZN(n1939)
         );
  BUF_X2 U1701 ( .I(rd_ptr[0]), .Z(n450) );
  NAND4_X1 U1702 ( .A1(n1944), .A2(n1943), .A3(n1942), .A4(n1941), .ZN(n1960)
         );
  NAND4_X1 U1703 ( .A1(n1924), .A2(n1923), .A3(n1922), .A4(n1921), .ZN(n1940)
         );
  BUF_X2 U1704 ( .I(rd_ptr[0]), .Z(n455) );
  BUF_X2 U1705 ( .I(rd_ptr[0]), .Z(n454) );
  BUF_X2 U1706 ( .I(rd_ptr[0]), .Z(n453) );
  BUF_X2 U1707 ( .I(rd_ptr[0]), .Z(n452) );
  BUF_X2 U1708 ( .I(rd_ptr[0]), .Z(n451) );
  INV_X1 U1709 ( .I(nxt_wr_ptr[0]), .ZN(n643) );
  MUX2_X1 U1710 ( .I0(queue[0]), .I1(queue[64]), .S(n455), .Z(N182) );
  MUX2_X1 U1711 ( .I0(queue[1]), .I1(queue[65]), .S(n455), .Z(N183) );
  MUX2_X1 U1712 ( .I0(queue[2]), .I1(queue[66]), .S(n455), .Z(N184) );
  MUX2_X1 U1713 ( .I0(queue[3]), .I1(queue[67]), .S(n455), .Z(N185) );
  MUX2_X1 U1714 ( .I0(queue[4]), .I1(queue[68]), .S(n455), .Z(N186) );
  MUX2_X1 U1715 ( .I0(queue[5]), .I1(queue[69]), .S(n455), .Z(N187) );
  MUX2_X1 U1716 ( .I0(queue[6]), .I1(queue[70]), .S(n455), .Z(N188) );
  MUX2_X1 U1717 ( .I0(queue[7]), .I1(queue[71]), .S(n455), .Z(N189) );
  MUX2_X1 U1718 ( .I0(queue[8]), .I1(queue[72]), .S(n455), .Z(N190) );
  MUX2_X1 U1719 ( .I0(queue[9]), .I1(queue[73]), .S(n455), .Z(N191) );
  MUX2_X1 U1720 ( .I0(queue[10]), .I1(queue[74]), .S(n455), .Z(N192) );
  MUX2_X1 U1721 ( .I0(queue[11]), .I1(queue[75]), .S(n455), .Z(N193) );
  MUX2_X1 U1722 ( .I0(queue[12]), .I1(queue[76]), .S(n454), .Z(N194) );
  MUX2_X1 U1723 ( .I0(queue[13]), .I1(queue[77]), .S(n454), .Z(N195) );
  MUX2_X1 U1724 ( .I0(queue[14]), .I1(queue[78]), .S(n454), .Z(N196) );
  MUX2_X1 U1725 ( .I0(queue[15]), .I1(queue[79]), .S(n454), .Z(N197) );
  MUX2_X1 U1726 ( .I0(queue[16]), .I1(queue[80]), .S(n454), .Z(N198) );
  MUX2_X1 U1727 ( .I0(queue[17]), .I1(queue[81]), .S(n454), .Z(N199) );
  MUX2_X1 U1728 ( .I0(queue[18]), .I1(queue[82]), .S(n454), .Z(N200) );
  MUX2_X1 U1729 ( .I0(queue[19]), .I1(queue[83]), .S(n454), .Z(N201) );
  MUX2_X1 U1730 ( .I0(queue[20]), .I1(queue[84]), .S(n454), .Z(N202) );
  MUX2_X1 U1731 ( .I0(queue[21]), .I1(queue[85]), .S(n454), .Z(N203) );
  MUX2_X1 U1732 ( .I0(queue[22]), .I1(queue[86]), .S(n454), .Z(N204) );
  MUX2_X1 U1733 ( .I0(queue[23]), .I1(queue[87]), .S(n454), .Z(N205) );
  MUX2_X1 U1734 ( .I0(queue[24]), .I1(queue[88]), .S(n453), .Z(N206) );
  MUX2_X1 U1735 ( .I0(queue[25]), .I1(queue[89]), .S(n453), .Z(N207) );
  MUX2_X1 U1736 ( .I0(queue[26]), .I1(queue[90]), .S(n453), .Z(N208) );
  MUX2_X1 U1737 ( .I0(queue[27]), .I1(queue[91]), .S(n453), .Z(N209) );
  MUX2_X1 U1738 ( .I0(queue[28]), .I1(queue[92]), .S(n453), .Z(N210) );
  MUX2_X1 U1739 ( .I0(queue[29]), .I1(queue[93]), .S(n453), .Z(N211) );
  MUX2_X1 U1740 ( .I0(queue[30]), .I1(queue[94]), .S(n453), .Z(N212) );
  MUX2_X1 U1741 ( .I0(queue[31]), .I1(queue[95]), .S(n453), .Z(N213) );
  MUX2_X1 U1742 ( .I0(queue[32]), .I1(queue[96]), .S(n453), .Z(N214) );
  MUX2_X1 U1743 ( .I0(queue[33]), .I1(queue[97]), .S(n453), .Z(N215) );
  MUX2_X1 U1744 ( .I0(queue[34]), .I1(queue[98]), .S(n453), .Z(N216) );
  MUX2_X1 U1745 ( .I0(queue[35]), .I1(queue[99]), .S(n453), .Z(N217) );
  MUX2_X1 U1746 ( .I0(queue[36]), .I1(queue[100]), .S(n452), .Z(N218) );
  MUX2_X1 U1747 ( .I0(queue[37]), .I1(queue[101]), .S(n452), .Z(N219) );
  MUX2_X1 U1748 ( .I0(queue[38]), .I1(queue[102]), .S(n452), .Z(N220) );
  MUX2_X1 U1749 ( .I0(queue[39]), .I1(queue[103]), .S(n452), .Z(N221) );
  MUX2_X1 U1750 ( .I0(queue[40]), .I1(queue[104]), .S(n452), .Z(N222) );
  MUX2_X1 U1751 ( .I0(queue[41]), .I1(queue[105]), .S(n452), .Z(N223) );
  MUX2_X1 U1752 ( .I0(queue[42]), .I1(queue[106]), .S(n452), .Z(N224) );
  MUX2_X1 U1753 ( .I0(queue[43]), .I1(queue[107]), .S(n452), .Z(N225) );
  MUX2_X1 U1754 ( .I0(queue[44]), .I1(queue[108]), .S(n452), .Z(N226) );
  MUX2_X1 U1755 ( .I0(queue[45]), .I1(queue[109]), .S(n452), .Z(N227) );
  MUX2_X1 U1756 ( .I0(queue[46]), .I1(queue[110]), .S(n452), .Z(N228) );
  MUX2_X1 U1757 ( .I0(queue[47]), .I1(queue[111]), .S(n452), .Z(N229) );
  MUX2_X1 U1758 ( .I0(queue[48]), .I1(queue[112]), .S(n451), .Z(N230) );
  MUX2_X1 U1759 ( .I0(queue[49]), .I1(queue[113]), .S(n451), .Z(N231) );
  MUX2_X1 U1760 ( .I0(queue[50]), .I1(queue[114]), .S(n451), .Z(N232) );
  MUX2_X1 U1761 ( .I0(queue[51]), .I1(queue[115]), .S(n451), .Z(N233) );
  MUX2_X1 U1762 ( .I0(queue[52]), .I1(queue[116]), .S(n451), .Z(N234) );
  MUX2_X1 U1763 ( .I0(queue[53]), .I1(queue[117]), .S(n451), .Z(N235) );
  MUX2_X1 U1764 ( .I0(queue[54]), .I1(queue[118]), .S(n451), .Z(N236) );
  MUX2_X1 U1765 ( .I0(queue[55]), .I1(queue[119]), .S(n451), .Z(N237) );
  MUX2_X1 U1766 ( .I0(queue[56]), .I1(queue[120]), .S(n451), .Z(N238) );
  MUX2_X1 U1767 ( .I0(queue[57]), .I1(queue[121]), .S(n451), .Z(N239) );
  MUX2_X1 U1768 ( .I0(queue[58]), .I1(queue[122]), .S(n451), .Z(N240) );
  MUX2_X1 U1769 ( .I0(queue[59]), .I1(queue[123]), .S(n451), .Z(N241) );
  MUX2_X1 U1770 ( .I0(queue[60]), .I1(queue[124]), .S(n450), .Z(N242) );
  MUX2_X1 U1771 ( .I0(queue[61]), .I1(queue[125]), .S(n450), .Z(N243) );
  MUX2_X1 U1772 ( .I0(queue[62]), .I1(queue[126]), .S(n450), .Z(N244) );
  MUX2_X1 U1773 ( .I0(queue[63]), .I1(queue[127]), .S(n450), .Z(N245) );
  INV_X1 U1774 ( .I(n565), .ZN(n537) );
  INV_X1 U1775 ( .I(n525), .ZN(n538) );
  INV_X1 U1776 ( .I(n525), .ZN(n539) );
  INV_X1 U1777 ( .I(n525), .ZN(n540) );
  INV_X1 U1778 ( .I(n526), .ZN(n541) );
  INV_X1 U1779 ( .I(n526), .ZN(n542) );
  INV_X1 U1780 ( .I(n526), .ZN(n543) );
  INV_X1 U1781 ( .I(n527), .ZN(n544) );
  INV_X1 U1782 ( .I(n527), .ZN(n545) );
  INV_X1 U1783 ( .I(n527), .ZN(n546) );
  INV_X1 U1784 ( .I(n527), .ZN(n547) );
  INV_X1 U1785 ( .I(n528), .ZN(n548) );
  INV_X1 U1786 ( .I(n528), .ZN(n549) );
  INV_X1 U1787 ( .I(n528), .ZN(n550) );
  INV_X1 U1788 ( .I(n528), .ZN(n551) );
  INV_X1 U1789 ( .I(n528), .ZN(n552) );
  INV_X1 U1790 ( .I(n529), .ZN(n553) );
  INV_X1 U1791 ( .I(n529), .ZN(n554) );
  INV_X1 U1792 ( .I(n529), .ZN(n555) );
  INV_X1 U1793 ( .I(n529), .ZN(n556) );
  INV_X1 U1794 ( .I(n529), .ZN(n557) );
  INV_X1 U1795 ( .I(n530), .ZN(n558) );
  INV_X1 U1796 ( .I(n530), .ZN(n559) );
  INV_X1 U1797 ( .I(n530), .ZN(n560) );
  INV_X1 U1798 ( .I(n530), .ZN(n561) );
  INV_X1 U1799 ( .I(n530), .ZN(n562) );
  INV_X1 U1800 ( .I(n531), .ZN(n563) );
  INV_X1 U1801 ( .I(n531), .ZN(n564) );
  INV_X1 U1802 ( .I(n531), .ZN(n565) );
endmodule


module pe_front_end_GENE_SZ64_ATTR_SZ8 ( clk, rst, bubble, bias, gene1_in, 
        gene2_in, gene1_out, gene2_out );
  input [63:0] gene1_in;
  input [63:0] gene2_in;
  output [63:0] gene1_out;
  output [63:0] gene2_out;
  input clk, rst;
  output bubble, bias;
  wire   gene1_rd, gene2_rd, N2, N3, N6, N7, N142, N143, N144, N145, N146,
         N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157,
         N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168,
         N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179,
         N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190,
         N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201,
         N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212,
         N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223,
         N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234,
         N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245,
         N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256,
         N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267,
         N268, N269, N270, N271, N273, n143, n144, n145, n146, n1, n2, n3, n4,
         n5, n6, n139, n140, n141, n142, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212;
  wire   [63:0] gene1_q_out;
  wire   [63:0] gene2_q_out;

  DFFSNQ_X1 gene2_rd_reg ( .D(N142), .CLK(clk), .SN(1'b1), .Q(gene2_rd) );
  DFFSNQ_X1 gene1_rd_reg ( .D(n148), .CLK(clk), .SN(1'b1), .Q(gene1_rd) );
  DFFSNQ_X1 gene2_out_reg_46_ ( .D(N253), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[46]) );
  DFFSNQ_X1 gene2_out_reg_45_ ( .D(N252), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[45]) );
  DFFSNQ_X1 gene2_out_reg_44_ ( .D(N251), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[44]) );
  DFFSNQ_X1 gene2_out_reg_43_ ( .D(N250), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[43]) );
  DFFSNQ_X1 gene2_out_reg_42_ ( .D(N249), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[42]) );
  DFFSNQ_X1 gene2_out_reg_41_ ( .D(N248), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[41]) );
  DFFSNQ_X1 gene2_out_reg_40_ ( .D(N247), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[40]) );
  DFFSNQ_X1 gene2_out_reg_39_ ( .D(N246), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[39]) );
  DFFSNQ_X1 gene2_out_reg_38_ ( .D(N245), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[38]) );
  DFFSNQ_X1 gene2_out_reg_37_ ( .D(N244), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[37]) );
  DFFSNQ_X1 gene2_out_reg_36_ ( .D(N243), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[36]) );
  DFFSNQ_X1 gene2_out_reg_35_ ( .D(N242), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[35]) );
  DFFSNQ_X1 gene2_out_reg_34_ ( .D(N241), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[34]) );
  DFFSNQ_X1 gene2_out_reg_33_ ( .D(N240), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[33]) );
  DFFSNQ_X1 gene2_out_reg_32_ ( .D(N239), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[32]) );
  DFFSNQ_X1 gene2_out_reg_31_ ( .D(N238), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[31]) );
  DFFSNQ_X1 gene2_out_reg_30_ ( .D(N237), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[30]) );
  DFFSNQ_X1 gene2_out_reg_29_ ( .D(N236), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[29]) );
  DFFSNQ_X1 gene2_out_reg_28_ ( .D(N235), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[28]) );
  DFFSNQ_X1 gene2_out_reg_27_ ( .D(N234), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[27]) );
  DFFSNQ_X1 gene2_out_reg_26_ ( .D(N233), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[26]) );
  DFFSNQ_X1 gene2_out_reg_25_ ( .D(N232), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[25]) );
  DFFSNQ_X1 gene2_out_reg_24_ ( .D(N231), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[24]) );
  DFFSNQ_X1 gene2_out_reg_23_ ( .D(N230), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[23]) );
  DFFSNQ_X1 gene2_out_reg_22_ ( .D(N229), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[22]) );
  DFFSNQ_X1 gene2_out_reg_21_ ( .D(N228), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[21]) );
  DFFSNQ_X1 gene2_out_reg_20_ ( .D(N227), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[20]) );
  DFFSNQ_X1 gene2_out_reg_19_ ( .D(N226), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[19]) );
  DFFSNQ_X1 gene2_out_reg_18_ ( .D(N225), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[18]) );
  DFFSNQ_X1 gene2_out_reg_17_ ( .D(N224), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[17]) );
  DFFSNQ_X1 gene2_out_reg_16_ ( .D(N223), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[16]) );
  DFFSNQ_X1 gene2_out_reg_15_ ( .D(N222), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[15]) );
  DFFSNQ_X1 gene2_out_reg_14_ ( .D(N221), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[14]) );
  DFFSNQ_X1 gene2_out_reg_13_ ( .D(N220), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[13]) );
  DFFSNQ_X1 gene2_out_reg_12_ ( .D(N219), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[12]) );
  DFFSNQ_X1 gene2_out_reg_11_ ( .D(N218), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[11]) );
  DFFSNQ_X1 gene2_out_reg_10_ ( .D(N217), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[10]) );
  DFFSNQ_X1 gene2_out_reg_9_ ( .D(N216), .CLK(clk), .SN(1'b1), .Q(gene2_out[9]) );
  DFFSNQ_X1 gene2_out_reg_8_ ( .D(N215), .CLK(clk), .SN(1'b1), .Q(gene2_out[8]) );
  DFFSNQ_X1 gene2_out_reg_7_ ( .D(N214), .CLK(clk), .SN(1'b1), .Q(gene2_out[7]) );
  DFFSNQ_X1 gene2_out_reg_6_ ( .D(N213), .CLK(clk), .SN(1'b1), .Q(gene2_out[6]) );
  DFFSNQ_X1 gene2_out_reg_5_ ( .D(N212), .CLK(clk), .SN(1'b1), .Q(gene2_out[5]) );
  DFFSNQ_X1 gene2_out_reg_4_ ( .D(N211), .CLK(clk), .SN(1'b1), .Q(gene2_out[4]) );
  DFFSNQ_X1 gene2_out_reg_3_ ( .D(N210), .CLK(clk), .SN(1'b1), .Q(gene2_out[3]) );
  DFFSNQ_X1 gene2_out_reg_2_ ( .D(N209), .CLK(clk), .SN(1'b1), .Q(gene2_out[2]) );
  DFFSNQ_X1 gene2_out_reg_1_ ( .D(N208), .CLK(clk), .SN(1'b1), .Q(gene2_out[1]) );
  DFFSNQ_X1 gene2_out_reg_0_ ( .D(N207), .CLK(clk), .SN(1'b1), .Q(gene2_out[0]) );
  DFFSNQ_X1 gene1_out_reg_0_ ( .D(N143), .CLK(clk), .SN(1'b1), .Q(gene1_out[0]) );
  DFFSNQ_X1 gene1_out_reg_1_ ( .D(N144), .CLK(clk), .SN(1'b1), .Q(gene1_out[1]) );
  DFFSNQ_X1 gene1_out_reg_2_ ( .D(N145), .CLK(clk), .SN(1'b1), .Q(gene1_out[2]) );
  DFFSNQ_X1 gene1_out_reg_3_ ( .D(N146), .CLK(clk), .SN(1'b1), .Q(gene1_out[3]) );
  DFFSNQ_X1 gene1_out_reg_4_ ( .D(N147), .CLK(clk), .SN(1'b1), .Q(gene1_out[4]) );
  DFFSNQ_X1 gene1_out_reg_5_ ( .D(N148), .CLK(clk), .SN(1'b1), .Q(gene1_out[5]) );
  DFFSNQ_X1 gene1_out_reg_6_ ( .D(N149), .CLK(clk), .SN(1'b1), .Q(gene1_out[6]) );
  DFFSNQ_X1 gene1_out_reg_7_ ( .D(N150), .CLK(clk), .SN(1'b1), .Q(gene1_out[7]) );
  DFFSNQ_X1 gene1_out_reg_8_ ( .D(N151), .CLK(clk), .SN(1'b1), .Q(gene1_out[8]) );
  DFFSNQ_X1 gene1_out_reg_9_ ( .D(N152), .CLK(clk), .SN(1'b1), .Q(gene1_out[9]) );
  DFFSNQ_X1 gene1_out_reg_10_ ( .D(N153), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[10]) );
  DFFSNQ_X1 gene1_out_reg_11_ ( .D(N154), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[11]) );
  DFFSNQ_X1 gene1_out_reg_12_ ( .D(N155), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[12]) );
  DFFSNQ_X1 gene1_out_reg_13_ ( .D(N156), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[13]) );
  DFFSNQ_X1 gene1_out_reg_14_ ( .D(N157), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[14]) );
  DFFSNQ_X1 gene1_out_reg_15_ ( .D(N158), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[15]) );
  DFFSNQ_X1 gene1_out_reg_16_ ( .D(N159), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[16]) );
  DFFSNQ_X1 gene1_out_reg_17_ ( .D(N160), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[17]) );
  DFFSNQ_X1 gene1_out_reg_18_ ( .D(N161), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[18]) );
  DFFSNQ_X1 gene1_out_reg_19_ ( .D(N162), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[19]) );
  DFFSNQ_X1 gene1_out_reg_20_ ( .D(N163), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[20]) );
  DFFSNQ_X1 gene1_out_reg_21_ ( .D(N164), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[21]) );
  DFFSNQ_X1 gene1_out_reg_22_ ( .D(N165), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[22]) );
  DFFSNQ_X1 gene1_out_reg_23_ ( .D(N166), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[23]) );
  DFFSNQ_X1 gene1_out_reg_24_ ( .D(N167), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[24]) );
  DFFSNQ_X1 gene1_out_reg_25_ ( .D(N168), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[25]) );
  DFFSNQ_X1 gene1_out_reg_26_ ( .D(N169), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[26]) );
  DFFSNQ_X1 gene1_out_reg_27_ ( .D(N170), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[27]) );
  DFFSNQ_X1 gene1_out_reg_28_ ( .D(N171), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[28]) );
  DFFSNQ_X1 gene1_out_reg_29_ ( .D(N172), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[29]) );
  DFFSNQ_X1 gene1_out_reg_30_ ( .D(N173), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[30]) );
  DFFSNQ_X1 gene1_out_reg_31_ ( .D(N174), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[31]) );
  DFFSNQ_X1 gene1_out_reg_32_ ( .D(N175), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[32]) );
  DFFSNQ_X1 gene1_out_reg_33_ ( .D(N176), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[33]) );
  DFFSNQ_X1 gene1_out_reg_34_ ( .D(N177), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[34]) );
  DFFSNQ_X1 gene1_out_reg_35_ ( .D(N178), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[35]) );
  DFFSNQ_X1 gene1_out_reg_36_ ( .D(N179), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[36]) );
  DFFSNQ_X1 gene1_out_reg_37_ ( .D(N180), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[37]) );
  DFFSNQ_X1 gene1_out_reg_38_ ( .D(N181), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[38]) );
  DFFSNQ_X1 gene1_out_reg_39_ ( .D(N182), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[39]) );
  DFFSNQ_X1 gene1_out_reg_40_ ( .D(N183), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[40]) );
  DFFSNQ_X1 gene1_out_reg_41_ ( .D(N184), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[41]) );
  DFFSNQ_X1 gene1_out_reg_42_ ( .D(N185), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[42]) );
  DFFSNQ_X1 gene1_out_reg_43_ ( .D(N186), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[43]) );
  DFFSNQ_X1 gene1_out_reg_44_ ( .D(N187), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[44]) );
  DFFSNQ_X1 gene1_out_reg_45_ ( .D(N188), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[45]) );
  DFFSNQ_X1 gene1_out_reg_46_ ( .D(N189), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[46]) );
  DFFSNQ_X1 gene1_out_reg_47_ ( .D(N190), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[47]) );
  DFFSNQ_X1 gene1_out_reg_48_ ( .D(N191), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[48]) );
  DFFSNQ_X1 gene1_out_reg_49_ ( .D(N192), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[49]) );
  DFFSNQ_X1 gene1_out_reg_50_ ( .D(N193), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[50]) );
  DFFSNQ_X1 gene1_out_reg_51_ ( .D(N194), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[51]) );
  DFFSNQ_X1 gene1_out_reg_52_ ( .D(N195), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[52]) );
  DFFSNQ_X1 gene1_out_reg_53_ ( .D(N196), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[53]) );
  DFFSNQ_X1 gene1_out_reg_54_ ( .D(N197), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[54]) );
  DFFSNQ_X1 gene1_out_reg_55_ ( .D(N198), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[55]) );
  DFFSNQ_X1 gene1_out_reg_56_ ( .D(N199), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[56]) );
  DFFSNQ_X1 gene1_out_reg_57_ ( .D(N200), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[57]) );
  DFFSNQ_X1 gene1_out_reg_58_ ( .D(N201), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[58]) );
  DFFSNQ_X1 gene1_out_reg_59_ ( .D(N202), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[59]) );
  DFFSNQ_X1 gene1_out_reg_60_ ( .D(N203), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[60]) );
  DFFSNQ_X1 gene1_out_reg_61_ ( .D(N204), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[61]) );
  DFFSNQ_X1 gene1_out_reg_62_ ( .D(N205), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[62]) );
  DFFSNQ_X1 gene1_out_reg_63_ ( .D(N206), .CLK(clk), .SN(1'b1), .Q(
        gene1_out[63]) );
  DFFSNQ_X1 bias_reg ( .D(n209), .CLK(clk), .SN(1'b1), .Q(bias) );
  DFFSNQ_X1 gene2_out_reg_47_ ( .D(N254), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[47]) );
  DFFSNQ_X1 gene2_out_reg_48_ ( .D(N255), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[48]) );
  DFFSNQ_X1 gene2_out_reg_49_ ( .D(N256), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[49]) );
  DFFSNQ_X1 gene2_out_reg_50_ ( .D(N257), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[50]) );
  DFFSNQ_X1 gene2_out_reg_51_ ( .D(N258), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[51]) );
  DFFSNQ_X1 gene2_out_reg_52_ ( .D(N259), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[52]) );
  DFFSNQ_X1 gene2_out_reg_53_ ( .D(N260), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[53]) );
  DFFSNQ_X1 gene2_out_reg_54_ ( .D(N261), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[54]) );
  DFFSNQ_X1 gene2_out_reg_55_ ( .D(N262), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[55]) );
  DFFSNQ_X1 gene2_out_reg_56_ ( .D(N263), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[56]) );
  DFFSNQ_X1 gene2_out_reg_57_ ( .D(N264), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[57]) );
  DFFSNQ_X1 gene2_out_reg_58_ ( .D(N265), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[58]) );
  DFFSNQ_X1 gene2_out_reg_59_ ( .D(N266), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[59]) );
  DFFSNQ_X1 gene2_out_reg_60_ ( .D(N267), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[60]) );
  DFFSNQ_X1 gene2_out_reg_61_ ( .D(N268), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[61]) );
  DFFSNQ_X1 gene2_out_reg_62_ ( .D(N269), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[62]) );
  DFFSNQ_X1 gene2_out_reg_63_ ( .D(N270), .CLK(clk), .SN(1'b1), .Q(
        gene2_out[63]) );
  DFFSNQ_X1 bubble_reg ( .D(N271), .CLK(clk), .SN(1'b1), .Q(bubble) );
  AND2_X1 U147 ( .A1(gene2_q_out[63]), .A2(n1), .Z(N270) );
  AND2_X1 U148 ( .A1(gene2_q_out[62]), .A2(n1), .Z(N269) );
  AND2_X1 U149 ( .A1(gene2_q_out[61]), .A2(n1), .Z(N268) );
  AND2_X1 U150 ( .A1(gene2_q_out[60]), .A2(n1), .Z(N267) );
  AND2_X1 U151 ( .A1(gene2_q_out[59]), .A2(n1), .Z(N266) );
  AND2_X1 U152 ( .A1(gene2_q_out[58]), .A2(n1), .Z(N265) );
  AND2_X1 U153 ( .A1(gene2_q_out[57]), .A2(n1), .Z(N264) );
  AND2_X1 U154 ( .A1(gene2_q_out[56]), .A2(n1), .Z(N263) );
  AND2_X1 U155 ( .A1(gene2_q_out[55]), .A2(n1), .Z(N262) );
  AND2_X1 U156 ( .A1(gene2_q_out[54]), .A2(n1), .Z(N261) );
  AND2_X1 U157 ( .A1(gene2_q_out[53]), .A2(n1), .Z(N260) );
  AND2_X1 U158 ( .A1(gene2_q_out[52]), .A2(n1), .Z(N259) );
  AND2_X1 U159 ( .A1(gene2_q_out[51]), .A2(n2), .Z(N258) );
  AND2_X1 U160 ( .A1(gene2_q_out[50]), .A2(n2), .Z(N257) );
  AND2_X1 U161 ( .A1(gene2_q_out[49]), .A2(n2), .Z(N256) );
  AND2_X1 U162 ( .A1(gene2_q_out[48]), .A2(n2), .Z(N255) );
  AND2_X1 U163 ( .A1(gene2_q_out[47]), .A2(n2), .Z(N254) );
  AND2_X1 U164 ( .A1(gene2_q_out[46]), .A2(n2), .Z(N253) );
  AND2_X1 U165 ( .A1(gene2_q_out[45]), .A2(n2), .Z(N252) );
  AND2_X1 U166 ( .A1(gene2_q_out[44]), .A2(n2), .Z(N251) );
  AND2_X1 U167 ( .A1(gene2_q_out[43]), .A2(n2), .Z(N250) );
  AND2_X1 U168 ( .A1(gene2_q_out[42]), .A2(n2), .Z(N249) );
  AND2_X1 U169 ( .A1(gene2_q_out[41]), .A2(n2), .Z(N248) );
  AND2_X1 U170 ( .A1(gene2_q_out[40]), .A2(n2), .Z(N247) );
  AND2_X1 U171 ( .A1(gene2_q_out[39]), .A2(n3), .Z(N246) );
  AND2_X1 U172 ( .A1(gene2_q_out[38]), .A2(n3), .Z(N245) );
  AND2_X1 U173 ( .A1(gene2_q_out[37]), .A2(n3), .Z(N244) );
  AND2_X1 U174 ( .A1(gene2_q_out[36]), .A2(n3), .Z(N243) );
  AND2_X1 U175 ( .A1(gene2_q_out[35]), .A2(n3), .Z(N242) );
  AND2_X1 U176 ( .A1(gene2_q_out[34]), .A2(n3), .Z(N241) );
  AND2_X1 U177 ( .A1(gene2_q_out[33]), .A2(n3), .Z(N240) );
  AND2_X1 U178 ( .A1(gene2_q_out[32]), .A2(n3), .Z(N239) );
  AND2_X1 U179 ( .A1(gene2_q_out[31]), .A2(n3), .Z(N238) );
  AND2_X1 U180 ( .A1(gene2_q_out[30]), .A2(n3), .Z(N237) );
  AND2_X1 U181 ( .A1(gene2_q_out[29]), .A2(n3), .Z(N236) );
  AND2_X1 U182 ( .A1(gene2_q_out[28]), .A2(n3), .Z(N235) );
  AND2_X1 U183 ( .A1(gene2_q_out[27]), .A2(n4), .Z(N234) );
  AND2_X1 U184 ( .A1(gene2_q_out[26]), .A2(n4), .Z(N233) );
  AND2_X1 U185 ( .A1(gene2_q_out[25]), .A2(n4), .Z(N232) );
  AND2_X1 U186 ( .A1(gene2_q_out[24]), .A2(n4), .Z(N231) );
  AND2_X1 U187 ( .A1(gene2_q_out[23]), .A2(n4), .Z(N230) );
  AND2_X1 U188 ( .A1(gene2_q_out[22]), .A2(n4), .Z(N229) );
  AND2_X1 U189 ( .A1(gene2_q_out[21]), .A2(n4), .Z(N228) );
  AND2_X1 U190 ( .A1(gene2_q_out[20]), .A2(n4), .Z(N227) );
  AND2_X1 U191 ( .A1(gene2_q_out[19]), .A2(n4), .Z(N226) );
  AND2_X1 U192 ( .A1(gene2_q_out[18]), .A2(n4), .Z(N225) );
  AND2_X1 U193 ( .A1(gene2_q_out[17]), .A2(n4), .Z(N224) );
  AND2_X1 U194 ( .A1(gene2_q_out[16]), .A2(n4), .Z(N223) );
  AND2_X1 U195 ( .A1(gene2_q_out[15]), .A2(n5), .Z(N222) );
  AND2_X1 U196 ( .A1(gene2_q_out[14]), .A2(n5), .Z(N221) );
  AND2_X1 U197 ( .A1(gene2_q_out[13]), .A2(n5), .Z(N220) );
  AND2_X1 U198 ( .A1(gene2_q_out[12]), .A2(n5), .Z(N219) );
  AND2_X1 U199 ( .A1(gene2_q_out[11]), .A2(n5), .Z(N218) );
  AND2_X1 U200 ( .A1(gene2_q_out[10]), .A2(n5), .Z(N217) );
  AND2_X1 U201 ( .A1(gene2_q_out[9]), .A2(n5), .Z(N216) );
  AND2_X1 U202 ( .A1(gene2_q_out[8]), .A2(n5), .Z(N215) );
  AND2_X1 U203 ( .A1(gene2_q_out[7]), .A2(n5), .Z(N214) );
  AND2_X1 U204 ( .A1(gene2_q_out[6]), .A2(n5), .Z(N213) );
  AND2_X1 U205 ( .A1(gene2_q_out[5]), .A2(n5), .Z(N212) );
  AND2_X1 U206 ( .A1(gene2_q_out[4]), .A2(n5), .Z(N211) );
  AND2_X1 U207 ( .A1(gene2_q_out[3]), .A2(n6), .Z(N210) );
  AND2_X1 U208 ( .A1(gene2_q_out[2]), .A2(n6), .Z(N209) );
  AND2_X1 U209 ( .A1(gene2_q_out[1]), .A2(n6), .Z(N208) );
  AND2_X1 U210 ( .A1(gene2_q_out[0]), .A2(n6), .Z(N207) );
  AND2_X1 U211 ( .A1(gene1_q_out[63]), .A2(n148), .Z(N206) );
  AND2_X1 U212 ( .A1(gene1_q_out[62]), .A2(n148), .Z(N205) );
  AND2_X1 U213 ( .A1(gene1_q_out[61]), .A2(n148), .Z(N204) );
  AND2_X1 U214 ( .A1(gene1_q_out[60]), .A2(n148), .Z(N203) );
  AND2_X1 U215 ( .A1(gene1_q_out[59]), .A2(n147), .Z(N202) );
  AND2_X1 U216 ( .A1(gene1_q_out[58]), .A2(n147), .Z(N201) );
  AND2_X1 U217 ( .A1(gene1_q_out[57]), .A2(n147), .Z(N200) );
  AND2_X1 U218 ( .A1(gene1_q_out[56]), .A2(n147), .Z(N199) );
  AND2_X1 U219 ( .A1(gene1_q_out[55]), .A2(n147), .Z(N198) );
  AND2_X1 U220 ( .A1(gene1_q_out[54]), .A2(n147), .Z(N197) );
  AND2_X1 U221 ( .A1(gene1_q_out[53]), .A2(n147), .Z(N196) );
  AND2_X1 U222 ( .A1(gene1_q_out[52]), .A2(n147), .Z(N195) );
  AND2_X1 U223 ( .A1(gene1_q_out[51]), .A2(n147), .Z(N194) );
  AND2_X1 U224 ( .A1(gene1_q_out[50]), .A2(n147), .Z(N193) );
  AND2_X1 U225 ( .A1(gene1_q_out[49]), .A2(n147), .Z(N192) );
  AND2_X1 U226 ( .A1(gene1_q_out[48]), .A2(n147), .Z(N191) );
  AND2_X1 U227 ( .A1(gene1_q_out[47]), .A2(n142), .Z(N190) );
  AND2_X1 U228 ( .A1(gene1_q_out[46]), .A2(n142), .Z(N189) );
  AND2_X1 U229 ( .A1(gene1_q_out[45]), .A2(n142), .Z(N188) );
  AND2_X1 U230 ( .A1(gene1_q_out[44]), .A2(n142), .Z(N187) );
  AND2_X1 U231 ( .A1(gene1_q_out[43]), .A2(n142), .Z(N186) );
  AND2_X1 U232 ( .A1(gene1_q_out[42]), .A2(n142), .Z(N185) );
  AND2_X1 U233 ( .A1(gene1_q_out[41]), .A2(n142), .Z(N184) );
  AND2_X1 U234 ( .A1(gene1_q_out[40]), .A2(n142), .Z(N183) );
  AND2_X1 U235 ( .A1(gene1_q_out[39]), .A2(n142), .Z(N182) );
  AND2_X1 U236 ( .A1(gene1_q_out[38]), .A2(n142), .Z(N181) );
  AND2_X1 U237 ( .A1(gene1_q_out[37]), .A2(n142), .Z(N180) );
  AND2_X1 U238 ( .A1(gene1_q_out[36]), .A2(n142), .Z(N179) );
  AND2_X1 U239 ( .A1(gene1_q_out[35]), .A2(n141), .Z(N178) );
  AND2_X1 U240 ( .A1(gene1_q_out[34]), .A2(n141), .Z(N177) );
  AND2_X1 U241 ( .A1(gene1_q_out[33]), .A2(n141), .Z(N176) );
  AND2_X1 U242 ( .A1(gene1_q_out[32]), .A2(n141), .Z(N175) );
  AND2_X1 U243 ( .A1(gene1_q_out[31]), .A2(n141), .Z(N174) );
  AND2_X1 U244 ( .A1(gene1_q_out[30]), .A2(n141), .Z(N173) );
  AND2_X1 U245 ( .A1(gene1_q_out[29]), .A2(n141), .Z(N172) );
  AND2_X1 U246 ( .A1(gene1_q_out[28]), .A2(n141), .Z(N171) );
  AND2_X1 U247 ( .A1(gene1_q_out[27]), .A2(n141), .Z(N170) );
  AND2_X1 U248 ( .A1(gene1_q_out[26]), .A2(n141), .Z(N169) );
  AND2_X1 U249 ( .A1(gene1_q_out[25]), .A2(n141), .Z(N168) );
  AND2_X1 U250 ( .A1(gene1_q_out[24]), .A2(n141), .Z(N167) );
  AND2_X1 U251 ( .A1(gene1_q_out[23]), .A2(n140), .Z(N166) );
  AND2_X1 U252 ( .A1(gene1_q_out[22]), .A2(n140), .Z(N165) );
  AND2_X1 U253 ( .A1(gene1_q_out[21]), .A2(n140), .Z(N164) );
  AND2_X1 U254 ( .A1(gene1_q_out[20]), .A2(n140), .Z(N163) );
  AND2_X1 U255 ( .A1(gene1_q_out[19]), .A2(n140), .Z(N162) );
  AND2_X1 U256 ( .A1(gene1_q_out[18]), .A2(n140), .Z(N161) );
  AND2_X1 U257 ( .A1(gene1_q_out[17]), .A2(n140), .Z(N160) );
  AND2_X1 U258 ( .A1(gene1_q_out[16]), .A2(n140), .Z(N159) );
  AND2_X1 U259 ( .A1(gene1_q_out[15]), .A2(n140), .Z(N158) );
  AND2_X1 U260 ( .A1(gene1_q_out[14]), .A2(n140), .Z(N157) );
  AND2_X1 U261 ( .A1(gene1_q_out[13]), .A2(n140), .Z(N156) );
  AND2_X1 U262 ( .A1(gene1_q_out[12]), .A2(n140), .Z(N155) );
  AND2_X1 U263 ( .A1(gene1_q_out[11]), .A2(n139), .Z(N154) );
  AND2_X1 U264 ( .A1(gene1_q_out[10]), .A2(n139), .Z(N153) );
  AND2_X1 U265 ( .A1(gene1_q_out[9]), .A2(n139), .Z(N152) );
  AND2_X1 U266 ( .A1(gene1_q_out[8]), .A2(n139), .Z(N151) );
  AND2_X1 U267 ( .A1(gene1_q_out[7]), .A2(n139), .Z(N150) );
  AND2_X1 U268 ( .A1(gene1_q_out[6]), .A2(n139), .Z(N149) );
  AND2_X1 U269 ( .A1(gene1_q_out[5]), .A2(n139), .Z(N148) );
  AND2_X1 U270 ( .A1(gene1_q_out[4]), .A2(n139), .Z(N147) );
  AND2_X1 U271 ( .A1(gene1_q_out[3]), .A2(n139), .Z(N146) );
  AND2_X1 U272 ( .A1(gene1_q_out[2]), .A2(n139), .Z(N145) );
  AND2_X1 U273 ( .A1(gene1_q_out[1]), .A2(n139), .Z(N144) );
  AND2_X1 U274 ( .A1(gene1_q_out[0]), .A2(n139), .Z(N143) );
  OR2_X1 U275 ( .A1(n6), .A2(n209), .Z(N273) );
  circ_q_WORD_SZ64_1 gene1_q ( .clk(clk), .rst(rst), .rd(gene1_rd), .wr(1'b1), 
        .data_in(gene1_in), .data_out(gene1_q_out) );
  circ_q_WORD_SZ64_0 gene2_q ( .clk(clk), .rst(rst), .rd(gene2_rd), .wr(1'b1), 
        .data_in(gene2_in), .data_out(gene2_q_out) );
  BUF_X2 U4 ( .I(n144), .Z(n6) );
  BUF_X2 U5 ( .I(n144), .Z(n1) );
  BUF_X2 U137 ( .I(n144), .Z(n5) );
  BUF_X2 U138 ( .I(n144), .Z(n4) );
  BUF_X2 U139 ( .I(n144), .Z(n3) );
  BUF_X2 U140 ( .I(n144), .Z(n2) );
  NOR2_X1 U141 ( .A1(n212), .A2(n210), .ZN(n144) );
  BUF_X2 U142 ( .I(N273), .Z(n141) );
  BUF_X2 U143 ( .I(N273), .Z(n140) );
  BUF_X2 U144 ( .I(N273), .Z(n139) );
  BUF_X2 U145 ( .I(N273), .Z(n147) );
  BUF_X2 U146 ( .I(N273), .Z(n142) );
  BUF_X2 U276 ( .I(N273), .Z(n148) );
  INV_X1 U277 ( .I(N2), .ZN(n210) );
  INV_X1 U278 ( .I(N6), .ZN(n212) );
  NOR2_X1 U279 ( .A1(n211), .A2(N6), .ZN(n146) );
  INV_X1 U280 ( .I(n155), .ZN(n175) );
  INV_X1 U281 ( .I(n145), .ZN(n209) );
  AOI22_X1 U282 ( .A1(n210), .A2(N3), .B1(N2), .B2(n146), .ZN(n145) );
  INV_X1 U283 ( .I(n185), .ZN(n205) );
  OAI22_X1 U284 ( .A1(N3), .A2(N2), .B1(n210), .B2(n143), .ZN(N271) );
  NAND2_X1 U285 ( .A1(n212), .A2(n211), .ZN(n143) );
  OAI22_X1 U286 ( .A1(N3), .A2(N2), .B1(n146), .B2(n210), .ZN(N142) );
  INV_X1 U287 ( .I(N7), .ZN(n211) );
  INV_X1 U288 ( .I(gene2_q_out[40]), .ZN(n173) );
  INV_X1 U289 ( .I(gene1_q_out[42]), .ZN(n170) );
  INV_X1 U290 ( .I(gene2_q_out[41]), .ZN(n174) );
  INV_X1 U291 ( .I(gene2_q_out[43]), .ZN(n176) );
  INV_X1 U292 ( .I(gene1_q_out[44]), .ZN(n171) );
  INV_X1 U293 ( .I(gene2_q_out[32]), .ZN(n203) );
  INV_X1 U294 ( .I(gene1_q_out[34]), .ZN(n200) );
  INV_X1 U295 ( .I(gene1_q_out[46]), .ZN(n172) );
  INV_X1 U296 ( .I(gene2_q_out[45]), .ZN(n177) );
  INV_X1 U297 ( .I(gene2_q_out[33]), .ZN(n204) );
  INV_X1 U298 ( .I(gene2_q_out[47]), .ZN(n178) );
  INV_X1 U299 ( .I(gene2_q_out[35]), .ZN(n206) );
  INV_X1 U300 ( .I(gene1_q_out[36]), .ZN(n201) );
  INV_X1 U301 ( .I(gene1_q_out[38]), .ZN(n202) );
  INV_X1 U302 ( .I(gene2_q_out[37]), .ZN(n207) );
  INV_X1 U303 ( .I(gene2_q_out[39]), .ZN(n208) );
  AND2_X1 U304 ( .A1(gene1_q_out[40]), .A2(n173), .Z(n149) );
  OAI22_X1 U305 ( .A1(gene1_q_out[41]), .A2(n149), .B1(n149), .B2(n174), .ZN(
        n150) );
  OR2_X1 U306 ( .A1(n172), .A2(gene2_q_out[46]), .Z(n151) );
  NAND2_X1 U307 ( .A1(gene1_q_out[45]), .A2(n177), .ZN(n152) );
  OR2_X1 U308 ( .A1(n171), .A2(gene2_q_out[44]), .Z(n153) );
  NAND4_X1 U309 ( .A1(n150), .A2(n151), .A3(n152), .A4(n153), .ZN(n169) );
  NAND2_X1 U310 ( .A1(gene1_q_out[43]), .A2(n176), .ZN(n154) );
  NOR2_X1 U311 ( .A1(n170), .A2(gene2_q_out[42]), .ZN(n155) );
  NAND2_X1 U312 ( .A1(n154), .A2(n175), .ZN(n168) );
  AND2_X1 U313 ( .A1(gene1_q_out[47]), .A2(n178), .Z(n167) );
  AND2_X1 U314 ( .A1(n152), .A2(n151), .Z(n165) );
  AND2_X1 U315 ( .A1(n154), .A2(n153), .Z(n162) );
  OR2_X1 U316 ( .A1(n173), .A2(gene1_q_out[40]), .Z(n157) );
  OR2_X1 U317 ( .A1(n157), .A2(gene1_q_out[41]), .Z(n156) );
  AOI21_X1 U318 ( .A1(n156), .A2(n174), .B(n155), .ZN(n159) );
  NAND2_X1 U319 ( .A1(gene1_q_out[41]), .A2(n157), .ZN(n158) );
  AOI22_X1 U320 ( .A1(gene2_q_out[42]), .A2(n170), .B1(n159), .B2(n158), .ZN(
        n160) );
  OAI21_X1 U321 ( .A1(gene1_q_out[43]), .A2(n176), .B(n160), .ZN(n161) );
  AOI22_X1 U322 ( .A1(gene2_q_out[44]), .A2(n171), .B1(n162), .B2(n161), .ZN(
        n163) );
  OAI21_X1 U323 ( .A1(gene1_q_out[45]), .A2(n177), .B(n163), .ZN(n164) );
  AOI22_X1 U324 ( .A1(gene2_q_out[46]), .A2(n172), .B1(n165), .B2(n164), .ZN(
        n166) );
  OAI22_X1 U325 ( .A1(gene1_q_out[47]), .A2(n178), .B1(n167), .B2(n166), .ZN(
        N3) );
  NOR4_X1 U326 ( .A1(n169), .A2(n168), .A3(N3), .A4(n167), .ZN(N2) );
  AND2_X1 U327 ( .A1(gene1_q_out[32]), .A2(n203), .Z(n179) );
  OAI22_X1 U328 ( .A1(gene1_q_out[33]), .A2(n179), .B1(n179), .B2(n204), .ZN(
        n180) );
  OR2_X1 U329 ( .A1(n202), .A2(gene2_q_out[38]), .Z(n181) );
  NAND2_X1 U330 ( .A1(gene1_q_out[37]), .A2(n207), .ZN(n182) );
  OR2_X1 U331 ( .A1(n201), .A2(gene2_q_out[36]), .Z(n183) );
  NAND4_X1 U332 ( .A1(n180), .A2(n181), .A3(n182), .A4(n183), .ZN(n199) );
  NAND2_X1 U333 ( .A1(gene1_q_out[35]), .A2(n206), .ZN(n184) );
  NOR2_X1 U334 ( .A1(n200), .A2(gene2_q_out[34]), .ZN(n185) );
  NAND2_X1 U335 ( .A1(n184), .A2(n205), .ZN(n198) );
  AND2_X1 U336 ( .A1(gene1_q_out[39]), .A2(n208), .Z(n197) );
  AND2_X1 U337 ( .A1(n182), .A2(n181), .Z(n195) );
  AND2_X1 U338 ( .A1(n184), .A2(n183), .Z(n192) );
  OR2_X1 U339 ( .A1(n203), .A2(gene1_q_out[32]), .Z(n187) );
  OR2_X1 U340 ( .A1(n187), .A2(gene1_q_out[33]), .Z(n186) );
  AOI21_X1 U341 ( .A1(n186), .A2(n204), .B(n185), .ZN(n189) );
  NAND2_X1 U342 ( .A1(gene1_q_out[33]), .A2(n187), .ZN(n188) );
  AOI22_X1 U343 ( .A1(gene2_q_out[34]), .A2(n200), .B1(n189), .B2(n188), .ZN(
        n190) );
  OAI21_X1 U344 ( .A1(gene1_q_out[35]), .A2(n206), .B(n190), .ZN(n191) );
  AOI22_X1 U345 ( .A1(gene2_q_out[36]), .A2(n201), .B1(n192), .B2(n191), .ZN(
        n193) );
  OAI21_X1 U346 ( .A1(gene1_q_out[37]), .A2(n207), .B(n193), .ZN(n194) );
  AOI22_X1 U347 ( .A1(gene2_q_out[38]), .A2(n202), .B1(n195), .B2(n194), .ZN(
        n196) );
  OAI22_X1 U348 ( .A1(gene1_q_out[39]), .A2(n208), .B1(n197), .B2(n196), .ZN(
        N7) );
  NOR4_X1 U349 ( .A1(n199), .A2(n198), .A3(N7), .A4(n197), .ZN(N6) );
endmodule


module pe_front_end_wrapper ( clk, rst, gene_in1, gene_in2, clk_out );
  input [63:0] gene_in1;
  input [63:0] gene_in2;
  input clk, rst;
  output clk_out;
  wire   clk, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128;
  assign clk_out = clk;

  pe_front_end_GENE_SZ64_ATTR_SZ8 front_end ( .clk(clk), .rst(rst), .gene1_in(
        gene_in1), .gene2_in(gene_in2), .gene1_out({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64}), .gene2_out({SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128}) );
endmodule

